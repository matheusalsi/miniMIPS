#************************************************************************/
# Copyright        : (c) All Rights Reserved 
# Company          : X-FAB Semiconductor Foundries AG 
# Address          : Haarbergstr. 67,  D-99097 Erfurt, Germany 
#
# File             : D_CELLS.lef
# Description      : Layout Exchange Format
#                  
# Technology       : 018um
# Lib_version      : V 2.3.0
# Last Modified by : omy
# DATE             : Mar 30, 2011
# 
#************************************************************************/

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "<>" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE core
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.630 BY 4.880 ;
END core

MACRO SIGNALHOLD
    CLASS CORE ;
    FOREIGN SIGNALHOLD 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SIG
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.411  LAYER MET1  ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.260 1.730 1.600 2.080 ;
        RECT  0.730 1.640 1.320 2.020 ;
        RECT  0.980 1.240 1.320 2.020 ;
        RECT  0.180 1.785 1.600 2.020 ;
        RECT  0.180 2.895 0.520 3.235 ;
        RECT  0.180 1.785 0.420 3.235 ;
        END
    END SIG
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.980 -0.400 1.320 0.840 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.980 2.895 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.790 0.700 2.130 1.040 ;
        RECT  0.650 2.375 0.990 2.665 ;
        RECT  0.650 2.430 2.130 2.665 ;
        RECT  1.845 0.700 2.130 3.235 ;
        RECT  1.790 2.430 2.130 3.235 ;
    END
END SIGNALHOLD

MACRO SDFRX4
    CLASS CORE ;
    FOREIGN SDFRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.290  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.010 1.130 19.350 4.100 ;
        RECT  17.680 2.250 19.350 2.630 ;
        RECT  17.680 2.250 18.030 3.770 ;
        RECT  17.680 1.130 17.910 3.770 ;
        RECT  17.570 1.130 17.910 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.980 2.885 17.410 3.115 ;
        RECT  17.180 1.700 17.410 3.115 ;
        RECT  14.690 1.700 17.410 1.930 ;
        RECT  16.420 2.885 16.760 4.130 ;
        RECT  16.130 1.130 16.470 1.930 ;
        RECT  14.980 2.885 16.760 3.240 ;
        RECT  14.980 2.860 15.625 3.240 ;
        RECT  14.980 2.860 15.320 4.130 ;
        RECT  14.690 1.130 15.030 1.930 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.275 1.640 9.070 2.100 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.290 -0.400 18.630 1.470 ;
        RECT  16.850 -0.400 17.190 1.470 ;
        RECT  15.410 -0.400 15.750 1.470 ;
        RECT  13.095 -0.400 13.435 1.450 ;
        RECT  10.420 -0.400 10.760 1.370 ;
        RECT  8.415 -0.400 8.700 0.950 ;
        RECT  3.485 -0.400 4.935 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.250 4.170 18.590 5.280 ;
        RECT  17.130 4.170 17.470 5.280 ;
        RECT  15.700 3.470 16.040 5.280 ;
        RECT  14.220 4.160 14.560 5.280 ;
        RECT  12.960 3.510 13.300 5.280 ;
        RECT  10.940 3.965 11.280 5.280 ;
        RECT  8.545 2.910 8.830 5.280 ;
        RECT  4.475 3.965 4.815 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.960 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.400 5.335 1.740 ;
        RECT  3.895 1.400 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.070 1.190 6.395 1.530 ;
        RECT  5.620 1.300 6.395 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  5.620 1.300 5.850 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  5.620 2.935 6.045 3.275 ;
        RECT  4.630 3.045 6.045 3.275 ;
        RECT  6.425 2.980 6.765 3.735 ;
        RECT  2.020 3.505 6.765 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  5.165 0.630 6.855 0.860 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.165 0.630 5.395 1.170 ;
        RECT  2.255 0.940 5.395 1.170 ;
        RECT  6.625 0.630 6.855 1.660 ;
        RECT  6.625 1.320 7.210 1.660 ;
        RECT  8.930 0.775 10.190 1.005 ;
        RECT  7.085 0.735 7.955 1.090 ;
        RECT  7.595 0.735 7.955 1.410 ;
        RECT  8.930 0.775 9.160 1.410 ;
        RECT  7.595 1.180 9.160 1.410 ;
        RECT  9.960 0.775 10.190 1.960 ;
        RECT  9.960 1.730 11.670 1.960 ;
        RECT  11.330 1.730 11.670 2.070 ;
        RECT  7.595 0.735 7.855 2.940 ;
        RECT  12.000 1.540 12.340 1.880 ;
        RECT  6.080 1.840 6.390 2.195 ;
        RECT  6.080 1.965 7.365 2.195 ;
        RECT  9.390 1.240 9.730 2.680 ;
        RECT  9.390 2.340 10.310 2.680 ;
        RECT  12.000 1.540 12.230 2.680 ;
        RECT  8.085 2.450 12.230 2.680 ;
        RECT  7.025 1.965 7.365 3.400 ;
        RECT  8.085 2.450 8.315 3.400 ;
        RECT  7.025 3.170 8.315 3.400 ;
        RECT  9.210 2.450 9.520 3.855 ;
        RECT  10.410 3.505 11.750 3.735 ;
        RECT  11.520 3.505 11.750 4.100 ;
        RECT  9.210 3.625 10.640 3.855 ;
        RECT  11.520 3.760 12.030 4.100 ;
        RECT  11.570 0.970 11.910 1.310 ;
        RECT  11.570 1.080 12.800 1.310 ;
        RECT  13.460 2.355 13.800 2.700 ;
        RECT  12.570 2.470 13.800 2.700 ;
        RECT  12.570 1.080 12.800 3.220 ;
        RECT  9.750 2.990 12.800 3.220 ;
        RECT  11.930 2.990 12.270 3.330 ;
        RECT  9.750 2.990 10.090 3.395 ;
        RECT  13.940 1.070 14.280 1.910 ;
        RECT  13.030 1.680 14.280 1.910 ;
        RECT  13.030 1.680 13.370 2.030 ;
        RECT  14.050 2.310 16.950 2.540 ;
        RECT  16.610 2.310 16.950 2.650 ;
        RECT  14.050 1.070 14.280 3.160 ;
        RECT  13.660 2.930 14.280 3.160 ;
        RECT  13.660 2.930 14.000 3.760 ;
        RECT  1.145 1.585 2.80 1.815 ;
        RECT  2.020 3.505 5.80 3.735 ;
        RECT  2.255 0.940 4.70 1.170 ;
        RECT  8.085 2.450 11.00 2.680 ;
        RECT  9.750 2.990 11.60 3.220 ;
        RECT  14.050 2.310 15.50 2.540 ;
    END
END SDFRX4

MACRO SDFRX2
    CLASS CORE ;
    FOREIGN SDFRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.350 3.270 14.365 3.500 ;
        RECT  14.135 1.250 14.365 3.500 ;
        RECT  13.985 2.860 14.365 3.500 ;
        RECT  13.350 1.250 14.365 1.590 ;
        RECT  13.350 3.270 13.690 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.260 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.620 1.890 4.250 ;
        RECT  0.755 3.620 1.890 3.850 ;
        RECT  0.755 3.470 1.135 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.715 1.005 2.200 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.130 2.020 8.695 2.630 ;
        END
    END C
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 1.240 15.010 3.550 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.230 -0.400 15.570 0.720 ;
        RECT  14.110 -0.400 14.450 0.720 ;
        RECT  12.790 -0.400 13.130 0.720 ;
        RECT  11.385 -0.400 11.730 0.970 ;
        RECT  9.585 -0.400 9.925 0.790 ;
        RECT  7.560 -0.400 7.845 1.330 ;
        RECT  4.100 -0.400 4.440 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.230 3.950 15.570 5.280 ;
        RECT  14.110 3.950 14.450 5.280 ;
        RECT  12.590 4.125 12.930 5.280 ;
        RECT  11.185 3.960 11.525 5.280 ;
        RECT  9.005 3.660 9.345 5.280 ;
        RECT  7.705 3.530 8.045 5.280 ;
        RECT  4.415 4.100 4.755 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.160 2.015 ;
        RECT  4.890 1.785 5.160 2.485 ;
        RECT  3.480 1.400 3.710 3.240 ;
        RECT  3.480 2.900 4.200 3.240 ;
        RECT  5.330 1.205 5.670 1.545 ;
        RECT  3.940 2.245 4.660 2.585 ;
        RECT  4.430 2.245 4.660 2.945 ;
        RECT  4.430 2.715 5.620 2.945 ;
        RECT  5.390 1.205 5.620 3.385 ;
        RECT  5.390 3.045 5.985 3.385 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  4.690 0.745 6.470 0.975 ;
        RECT  1.770 0.940 4.920 1.170 ;
        RECT  6.130 0.745 6.470 1.595 ;
        RECT  6.405 3.530 6.745 3.870 ;
        RECT  2.120 3.640 6.745 3.870 ;
        RECT  2.120 3.640 2.410 4.020 ;
        RECT  8.075 0.680 9.355 0.910 ;
        RECT  6.785 0.630 7.125 0.965 ;
        RECT  9.125 0.680 9.355 1.250 ;
        RECT  9.125 1.020 9.615 1.250 ;
        RECT  9.385 1.020 9.615 1.920 ;
        RECT  8.075 0.680 8.305 1.790 ;
        RECT  6.895 1.560 8.305 1.790 ;
        RECT  9.385 1.690 10.550 1.920 ;
        RECT  10.210 1.690 10.550 2.030 ;
        RECT  6.895 0.630 7.125 2.165 ;
        RECT  6.520 1.825 7.285 2.165 ;
        RECT  6.945 1.560 7.285 2.825 ;
        RECT  8.535 1.140 8.895 1.710 ;
        RECT  8.535 1.480 9.155 1.710 ;
        RECT  5.850 1.900 6.190 2.625 ;
        RECT  5.850 2.395 6.445 2.625 ;
        RECT  9.675 2.360 11.060 2.700 ;
        RECT  8.925 2.470 11.060 2.700 ;
        RECT  7.515 2.020 7.800 3.300 ;
        RECT  6.215 2.395 6.445 3.300 ;
        RECT  7.515 2.960 9.155 3.300 ;
        RECT  8.925 1.480 9.155 3.300 ;
        RECT  6.215 3.055 9.155 3.300 ;
        RECT  10.560 0.630 10.900 0.970 ;
        RECT  10.670 0.630 10.900 1.460 ;
        RECT  10.670 1.230 11.520 1.460 ;
        RECT  11.290 1.230 11.520 3.160 ;
        RECT  12.370 2.750 12.655 3.160 ;
        RECT  10.155 2.930 12.655 3.160 ;
        RECT  10.155 2.930 10.495 3.825 ;
        RECT  12.090 0.680 12.430 2.520 ;
        RECT  11.750 2.290 13.380 2.520 ;
        RECT  11.750 2.290 12.040 2.650 ;
        RECT  12.885 2.290 13.380 2.650 ;
        RECT  12.885 2.290 13.115 3.720 ;
        RECT  12.030 3.390 13.115 3.720 ;
        RECT  1.770 0.940 3.60 1.170 ;
        RECT  2.120 3.640 5.60 3.870 ;
        RECT  8.925 2.470 10.30 2.700 ;
        RECT  6.215 3.055 8.20 3.300 ;
        RECT  10.155 2.930 11.40 3.160 ;
    END
END SDFRX2

MACRO SDFRX1
    CLASS CORE ;
    FOREIGN SDFRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.605 0.940 14.995 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 1.640 14.375 2.020 ;
        RECT  13.420 2.870 14.220 3.100 ;
        RECT  13.985 1.640 14.220 3.100 ;
        RECT  13.985 1.260 14.215 3.100 ;
        RECT  13.420 1.260 14.215 1.490 ;
        RECT  13.160 3.780 13.650 4.120 ;
        RECT  13.420 2.870 13.650 4.120 ;
        RECT  13.420 0.700 13.650 1.490 ;
        RECT  13.160 0.700 13.650 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 3.990 2.030 4.250 ;
        RECT  1.610 3.980 2.000 4.250 ;
        RECT  1.610 3.470 1.840 4.250 ;
        RECT  1.410 3.470 1.840 3.815 ;
        RECT  1.385 3.470 1.840 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.880 2.800 3.655 3.240 ;
        RECT  2.880 2.045 3.110 3.240 ;
        RECT  0.575 2.045 3.110 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 1.640 8.885 2.035 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.880 -0.400 14.220 1.030 ;
        RECT  12.000 -0.400 12.340 1.050 ;
        RECT  10.145 -0.400 10.485 1.030 ;
        RECT  8.085 -0.400 8.425 0.950 ;
        RECT  4.725 -0.400 5.065 0.655 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  2.825 1.090 3.825 1.320 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  13.880 3.330 14.220 5.280 ;
        RECT  12.365 4.040 12.705 5.280 ;
        RECT  9.480 3.500 9.820 5.280 ;
        RECT  8.180 3.620 8.520 5.280 ;
        RECT  4.905 3.845 5.230 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.630 1.815 ;
        RECT  3.290 1.555 3.630 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  3.900 1.755 4.240 2.110 ;
        RECT  3.900 1.880 5.275 2.110 ;
        RECT  4.935 1.880 5.275 2.220 ;
        RECT  3.900 1.755 4.215 3.425 ;
        RECT  5.885 1.200 6.225 1.540 ;
        RECT  4.445 2.565 4.775 3.155 ;
        RECT  5.680 1.310 5.920 3.155 ;
        RECT  4.445 2.925 6.460 3.155 ;
        RECT  6.120 2.925 6.460 3.460 ;
        RECT  2.255 0.630 4.495 0.860 ;
        RECT  5.295 0.630 7.025 0.860 ;
        RECT  4.265 0.630 4.495 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.295 0.630 5.525 1.115 ;
        RECT  4.265 0.885 5.525 1.115 ;
        RECT  6.685 0.630 7.025 1.685 ;
        RECT  2.070 3.420 2.410 3.760 ;
        RECT  4.445 3.385 5.710 3.615 ;
        RECT  5.480 3.385 5.710 3.930 ;
        RECT  2.070 3.530 3.580 3.760 ;
        RECT  4.445 3.385 4.675 3.885 ;
        RECT  3.365 3.655 4.675 3.885 ;
        RECT  6.880 3.620 7.220 3.930 ;
        RECT  5.480 3.700 7.220 3.930 ;
        RECT  9.115 1.095 9.455 1.460 ;
        RECT  6.165 2.165 6.505 2.675 ;
        RECT  7.745 2.105 8.095 2.460 ;
        RECT  6.165 2.445 7.010 2.675 ;
        RECT  9.115 1.095 9.345 3.120 ;
        RECT  8.940 2.890 10.730 3.120 ;
        RECT  6.780 2.445 7.010 3.390 ;
        RECT  7.990 2.245 8.220 3.390 ;
        RECT  8.940 2.710 9.170 3.390 ;
        RECT  10.390 2.890 10.730 3.230 ;
        RECT  6.780 3.160 9.170 3.390 ;
        RECT  8.655 0.630 9.915 0.860 ;
        RECT  7.285 0.645 7.625 1.410 ;
        RECT  8.655 0.630 8.885 1.410 ;
        RECT  7.285 1.180 8.885 1.410 ;
        RECT  6.965 1.915 7.515 2.205 ;
        RECT  9.685 0.630 9.915 2.450 ;
        RECT  9.685 2.220 10.465 2.450 ;
        RECT  10.125 2.330 11.210 2.560 ;
        RECT  7.285 0.645 7.515 2.930 ;
        RECT  7.285 2.690 7.760 2.930 ;
        RECT  10.980 2.330 11.210 3.320 ;
        RECT  10.980 2.980 11.405 3.320 ;
        RECT  10.995 0.710 11.670 1.070 ;
        RECT  11.440 2.430 11.885 2.660 ;
        RECT  11.440 0.710 11.670 2.660 ;
        RECT  11.650 2.660 12.520 3.000 ;
        RECT  11.650 2.430 11.880 3.840 ;
        RECT  10.630 3.550 11.880 3.840 ;
        RECT  11.900 1.615 13.195 1.955 ;
        RECT  12.960 1.615 13.195 2.475 ;
        RECT  11.900 1.615 12.185 2.135 ;
        RECT  12.960 2.135 13.355 2.475 ;
        RECT  12.960 1.615 13.190 3.470 ;
        RECT  12.460 3.240 13.190 3.470 ;
        RECT  12.460 3.240 12.800 3.580 ;
        RECT  1.255 1.585 2.80 1.815 ;
        RECT  4.445 2.925 5.40 3.155 ;
        RECT  2.255 0.630 3.90 0.860 ;
        RECT  6.780 3.160 8.50 3.390 ;
    END
END SDFRX1

MACRO SDFRX0
    CLASS CORE ;
    FOREIGN SDFRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.489  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.220 2.860 13.735 3.240 ;
        RECT  13.220 2.640 13.640 3.240 ;
        RECT  13.410 1.170 13.640 3.240 ;
        RECT  13.300 1.170 13.640 1.510 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.600  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 1.640 13.105 2.020 ;
        RECT  12.380 2.640 12.955 2.980 ;
        RECT  12.725 0.630 12.955 2.980 ;
        RECT  12.045 0.630 12.955 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.215 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.215 3.320 ;
        RECT  2.190 2.860 3.215 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.480 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.625 2.185 8.120 2.675 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  13.220 3.470 13.560 5.280 ;
        RECT  11.730 4.165 12.070 5.280 ;
        RECT  10.755 3.930 11.040 5.280 ;
        RECT  8.120 3.630 8.460 5.280 ;
        RECT  7.395 3.925 7.735 5.280 ;
        RECT  3.200 4.170 4.495 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.300 -0.400 13.640 0.710 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  9.270 -0.400 9.555 0.710 ;
        RECT  9.250 -0.400 9.555 0.675 ;
        RECT  7.375 -0.400 7.660 0.970 ;
        RECT  3.970 -0.400 4.310 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.215 1.815 ;
        RECT  2.930 1.585 3.215 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.445 1.805 4.770 2.035 ;
        RECT  3.445 1.805 3.875 2.095 ;
        RECT  3.445 1.805 3.835 2.105 ;
        RECT  4.485 1.805 4.770 2.205 ;
        RECT  3.445 1.805 3.675 3.425 ;
        RECT  3.445 3.085 4.195 3.425 ;
        RECT  5.000 1.230 5.800 1.540 ;
        RECT  3.905 2.325 4.190 2.665 ;
        RECT  3.905 2.435 5.230 2.665 ;
        RECT  5.000 1.230 5.230 3.480 ;
        RECT  4.995 2.435 5.230 3.480 ;
        RECT  4.995 3.250 5.725 3.480 ;
        RECT  5.385 3.250 5.725 3.790 ;
        RECT  4.540 0.640 6.500 0.920 ;
        RECT  6.160 0.640 6.500 0.980 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  4.540 0.640 4.770 1.355 ;
        RECT  1.980 1.125 4.770 1.355 ;
        RECT  1.995 3.710 5.050 3.940 ;
        RECT  4.820 3.710 5.050 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.185 3.925 6.525 4.250 ;
        RECT  4.820 4.020 6.525 4.250 ;
        RECT  5.460 2.440 5.800 2.780 ;
        RECT  7.045 2.355 7.395 2.695 ;
        RECT  5.460 2.530 6.190 2.780 ;
        RECT  8.350 2.600 9.410 2.940 ;
        RECT  8.350 1.230 8.580 3.245 ;
        RECT  7.165 2.905 8.580 3.245 ;
        RECT  5.960 2.530 6.190 3.695 ;
        RECT  7.165 2.355 7.395 3.695 ;
        RECT  5.960 3.465 7.395 3.695 ;
        RECT  7.890 0.770 9.040 1.000 ;
        RECT  7.890 0.770 8.120 1.480 ;
        RECT  6.865 1.250 8.120 1.480 ;
        RECT  8.810 0.770 9.040 2.160 ;
        RECT  6.865 1.250 7.205 2.110 ;
        RECT  5.460 1.770 7.205 2.110 ;
        RECT  8.810 1.930 9.635 2.160 ;
        RECT  9.295 2.040 9.955 2.270 ;
        RECT  6.585 1.770 6.815 3.230 ;
        RECT  6.585 2.895 6.930 3.230 ;
        RECT  9.725 2.040 9.955 3.400 ;
        RECT  6.585 2.900 6.935 3.230 ;
        RECT  9.725 3.060 10.065 3.400 ;
        RECT  10.125 1.110 10.525 1.450 ;
        RECT  11.390 2.340 11.680 2.680 ;
        RECT  10.295 2.450 11.680 2.680 ;
        RECT  10.295 1.110 10.525 3.970 ;
        RECT  9.350 3.630 10.525 3.970 ;
        RECT  12.045 1.350 12.385 2.320 ;
        RECT  11.085 1.670 12.385 2.010 ;
        RECT  11.910 1.980 12.495 2.320 ;
        RECT  11.910 1.670 12.140 3.335 ;
        RECT  11.130 3.105 12.140 3.335 ;
        RECT  11.130 3.105 11.470 3.445 ;
        RECT  0.980 1.585 2.60 1.815 ;
        RECT  1.980 1.125 3.80 1.355 ;
        RECT  1.995 3.710 4.50 3.940 ;
    END
END SDFRX0

MACRO SDFRSX4
    CLASS CORE ;
    FOREIGN SDFRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.085  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 1.130 19.980 3.060 ;
        RECT  18.360 2.250 19.980 2.630 ;
        RECT  18.360 2.250 18.715 3.060 ;
        RECT  18.360 1.130 18.590 3.060 ;
        RECT  18.200 1.130 18.590 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.090  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.635 2.880 18.065 3.110 ;
        RECT  17.835 1.700 18.065 3.110 ;
        RECT  15.535 1.700 18.065 1.930 ;
        RECT  15.635 2.880 17.415 3.240 ;
        RECT  16.760 1.130 17.100 1.930 ;
        RECT  15.635 2.860 16.255 3.240 ;
        RECT  15.635 2.860 15.975 4.100 ;
        RECT  15.535 0.700 15.765 1.930 ;
        RECT  15.280 0.700 15.765 1.040 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.760 1.640 14.365 2.070 ;
        END
    END SN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 1.660 9.500 2.100 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.470 ;
        RECT  17.480 -0.400 17.820 1.470 ;
        RECT  16.040 -0.400 16.380 1.470 ;
        RECT  13.480 -0.400 13.820 0.840 ;
        RECT  10.715 -0.400 11.000 1.370 ;
        RECT  8.820 -0.400 9.105 0.970 ;
        RECT  3.400 -0.400 5.150 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  19.000 3.295 19.340 5.280 ;
        RECT  17.705 3.555 18.045 5.280 ;
        RECT  16.355 3.470 16.695 5.280 ;
        RECT  14.875 4.140 15.215 5.280 ;
        RECT  13.590 2.890 13.930 5.280 ;
        RECT  11.370 3.965 11.710 5.280 ;
        RECT  8.975 2.910 9.260 5.280 ;
        RECT  4.795 3.965 5.135 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.585 5.740 1.875 ;
        RECT  5.400 1.585 5.740 2.265 ;
        RECT  3.895 1.585 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.475 1.190 6.800 1.530 ;
        RECT  6.025 1.300 6.800 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  6.025 1.300 6.255 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  6.025 2.935 6.450 3.275 ;
        RECT  4.630 3.045 6.450 3.275 ;
        RECT  6.830 2.980 7.170 3.735 ;
        RECT  2.020 3.505 7.170 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  5.380 0.630 7.260 0.860 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.380 0.630 5.610 1.170 ;
        RECT  2.255 0.940 5.610 1.170 ;
        RECT  7.030 0.630 7.260 1.660 ;
        RECT  7.030 1.320 7.615 1.660 ;
        RECT  9.335 0.775 10.485 1.005 ;
        RECT  7.490 0.735 8.360 1.090 ;
        RECT  8.000 0.735 8.360 1.430 ;
        RECT  9.335 0.775 9.565 1.430 ;
        RECT  8.000 1.200 9.565 1.430 ;
        RECT  10.255 0.775 10.485 1.960 ;
        RECT  10.255 1.730 11.910 1.960 ;
        RECT  11.570 1.730 11.910 2.070 ;
        RECT  8.000 0.735 8.285 2.940 ;
        RECT  6.485 1.840 6.795 2.195 ;
        RECT  6.485 1.965 7.770 2.195 ;
        RECT  9.795 1.240 10.025 2.680 ;
        RECT  9.795 2.340 10.740 2.680 ;
        RECT  12.240 1.540 12.525 2.680 ;
        RECT  8.515 2.450 12.525 2.680 ;
        RECT  9.640 2.450 9.980 2.860 ;
        RECT  7.430 1.965 7.770 3.400 ;
        RECT  8.515 2.450 8.745 3.400 ;
        RECT  7.430 3.170 8.745 3.400 ;
        RECT  9.640 2.450 9.870 3.855 ;
        RECT  10.840 3.505 12.180 3.735 ;
        RECT  11.950 3.505 12.180 4.100 ;
        RECT  9.640 3.625 11.070 3.855 ;
        RECT  11.950 3.760 12.460 4.100 ;
        RECT  11.810 0.970 12.150 1.310 ;
        RECT  11.810 1.080 12.985 1.310 ;
        RECT  14.505 2.320 14.845 2.660 ;
        RECT  12.755 2.430 14.845 2.660 ;
        RECT  12.755 1.080 12.985 3.220 ;
        RECT  10.180 2.990 12.985 3.220 ;
        RECT  12.360 2.990 12.700 3.330 ;
        RECT  10.180 2.990 10.520 3.395 ;
        RECT  13.215 1.180 15.050 1.410 ;
        RECT  14.710 1.180 15.050 1.700 ;
        RECT  13.215 1.180 13.500 1.530 ;
        RECT  14.710 1.470 15.305 1.700 ;
        RECT  15.075 2.310 17.605 2.540 ;
        RECT  17.265 2.310 17.605 2.650 ;
        RECT  15.075 1.470 15.305 3.120 ;
        RECT  14.315 2.890 15.305 3.120 ;
        RECT  14.315 2.890 14.655 3.730 ;
        RECT  1.145 1.585 2.70 1.815 ;
        RECT  2.020 3.505 6.70 3.735 ;
        RECT  2.255 0.940 4.30 1.170 ;
        RECT  8.515 2.450 11.20 2.680 ;
        RECT  12.755 2.430 13.60 2.660 ;
        RECT  10.180 2.990 11.80 3.220 ;
        RECT  15.075 2.310 16.90 2.540 ;
    END
END SDFRSX4

MACRO SDFRSX2
    CLASS CORE ;
    FOREIGN SDFRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.765 0.830 14.995 3.240 ;
        RECT  14.450 2.860 14.790 4.180 ;
        RECT  14.610 0.830 14.995 1.170 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.260 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.620 1.890 4.250 ;
        RECT  0.755 3.620 1.890 3.850 ;
        RECT  0.755 3.470 1.135 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.215 3.250 3.020 ;
        RECT  1.660 2.215 3.250 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.720 1.005 2.200 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 2.020 8.740 2.630 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.585 2.050 13.105 2.630 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.875 1.240 16.270 2.020 ;
        RECT  15.770 2.640 16.110 3.550 ;
        RECT  15.875 1.240 16.110 3.550 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 0.720 ;
        RECT  15.370 -0.400 15.710 0.720 ;
        RECT  13.850 -0.400 14.190 0.970 ;
        RECT  12.300 -0.400 12.645 1.090 ;
        RECT  9.910 -0.400 10.195 1.330 ;
        RECT  7.990 -0.400 8.275 1.330 ;
        RECT  4.530 -0.400 4.870 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.490 2.640 16.830 5.280 ;
        RECT  15.210 3.950 15.550 5.280 ;
        RECT  13.690 4.170 14.030 5.280 ;
        RECT  11.710 3.385 12.750 5.280 ;
        RECT  9.330 3.480 9.670 5.280 ;
        RECT  8.030 3.515 8.370 5.280 ;
        RECT  4.715 3.900 5.055 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.330 2.015 ;
        RECT  4.990 1.785 5.330 2.470 ;
        RECT  3.480 1.400 3.710 3.270 ;
        RECT  3.480 2.930 4.250 3.265 ;
        RECT  3.480 2.930 4.240 3.270 ;
        RECT  5.580 1.190 6.100 1.530 ;
        RECT  3.940 2.245 4.715 2.585 ;
        RECT  4.485 2.245 4.715 2.930 ;
        RECT  5.580 1.190 5.810 3.210 ;
        RECT  4.485 2.700 5.810 2.930 ;
        RECT  5.580 2.870 6.285 3.210 ;
        RECT  5.120 0.630 6.900 0.860 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  5.120 0.630 5.350 1.170 ;
        RECT  1.770 0.940 5.350 1.170 ;
        RECT  6.560 0.630 6.900 1.595 ;
        RECT  4.400 3.440 5.525 3.670 ;
        RECT  2.120 3.500 4.560 3.730 ;
        RECT  6.705 3.515 7.045 3.845 ;
        RECT  5.295 3.615 7.045 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  7.215 0.630 7.555 0.965 ;
        RECT  8.505 0.800 9.680 1.030 ;
        RECT  7.325 0.630 7.555 2.825 ;
        RECT  9.450 0.800 9.680 1.790 ;
        RECT  8.505 0.800 8.735 1.790 ;
        RECT  7.325 1.560 8.735 1.790 ;
        RECT  9.450 1.560 11.105 1.790 ;
        RECT  10.765 1.560 11.105 1.895 ;
        RECT  7.065 1.825 7.610 2.165 ;
        RECT  7.325 1.560 7.610 2.825 ;
        RECT  7.270 1.825 7.610 2.825 ;
        RECT  6.040 1.760 6.380 2.110 ;
        RECT  6.040 1.880 6.780 2.110 ;
        RECT  10.040 2.120 10.380 2.460 ;
        RECT  10.040 2.225 11.425 2.460 ;
        RECT  8.970 2.230 11.425 2.460 ;
        RECT  11.140 2.225 11.425 2.565 ;
        RECT  6.550 1.880 6.780 3.285 ;
        RECT  7.840 2.860 9.220 3.145 ;
        RECT  8.970 1.260 9.220 3.145 ;
        RECT  7.840 2.020 8.085 3.285 ;
        RECT  6.550 3.055 8.085 3.285 ;
        RECT  11.035 1.035 11.810 1.330 ;
        RECT  11.580 1.035 11.810 2.055 ;
        RECT  11.655 1.835 11.885 3.090 ;
        RECT  13.415 2.750 13.755 3.090 ;
        RECT  10.480 2.860 13.755 3.090 ;
        RECT  10.480 2.860 10.820 3.615 ;
        RECT  12.040 1.320 12.325 1.660 ;
        RECT  12.040 1.430 13.875 1.660 ;
        RECT  13.535 1.430 13.875 2.110 ;
        RECT  13.535 1.880 14.395 2.110 ;
        RECT  13.985 1.880 14.395 2.220 ;
        RECT  13.985 1.880 14.215 3.610 ;
        RECT  13.130 3.380 14.215 3.610 ;
        RECT  13.130 3.380 13.470 3.720 ;
        RECT  1.770 0.940 4.50 1.170 ;
        RECT  2.120 3.500 3.60 3.730 ;
        RECT  8.970 2.230 10.70 2.460 ;
        RECT  10.480 2.860 12.60 3.090 ;
    END
END SDFRSX2

MACRO SDFRSX1
    CLASS CORE ;
    FOREIGN SDFRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.855 1.640 9.375 2.110 ;
        END
    END C
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.850 2.860 16.255 3.240 ;
        RECT  15.850 0.940 16.190 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.165 1.640 15.620 2.020 ;
        RECT  14.520 2.870 15.395 3.100 ;
        RECT  15.165 1.235 15.395 3.100 ;
        RECT  14.570 1.235 15.395 1.465 ;
        RECT  14.570 0.700 14.800 1.465 ;
        RECT  14.410 3.625 14.750 3.965 ;
        RECT  14.520 2.870 14.750 3.965 ;
        RECT  14.410 0.700 14.800 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.670 3.995 2.030 4.250 ;
        RECT  1.670 3.960 2.015 4.250 ;
        RECT  1.670 3.470 1.900 4.250 ;
        RECT  1.410 3.470 1.900 3.815 ;
        RECT  1.385 3.470 1.900 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.940 2.800 3.655 3.190 ;
        RECT  2.940 2.045 3.170 3.190 ;
        RECT  0.575 2.045 3.170 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.805 2.710 3.190 ;
        RECT  2.370 2.505 2.710 3.190 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.075 2.250 13.735 2.700 ;
        END
    END SN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.130 -0.400 15.470 1.005 ;
        RECT  12.755 -0.400 13.095 1.025 ;
        RECT  10.770 -0.400 11.110 1.005 ;
        RECT  8.705 -0.400 9.045 0.950 ;
        RECT  5.170 -0.400 5.510 0.710 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  2.825 1.090 3.825 1.320 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.130 3.330 15.470 5.280 ;
        RECT  13.825 4.170 14.165 5.280 ;
        RECT  12.330 3.630 12.645 5.280 ;
        RECT  9.765 3.480 10.105 5.280 ;
        RECT  8.465 3.535 8.805 5.280 ;
        RECT  5.170 3.430 5.510 5.280 ;
        RECT  3.470 4.170 3.810 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.690 1.815 ;
        RECT  3.350 1.555 3.690 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  4.080 1.570 4.420 2.090 ;
        RECT  3.920 1.860 5.830 2.090 ;
        RECT  5.490 1.860 5.830 2.280 ;
        RECT  3.920 1.860 4.150 3.190 ;
        RECT  3.920 2.850 4.480 3.190 ;
        RECT  6.325 1.200 6.740 1.540 ;
        RECT  4.390 2.320 4.995 2.605 ;
        RECT  4.780 2.510 6.555 2.740 ;
        RECT  6.325 1.200 6.555 3.385 ;
        RECT  6.325 3.045 6.745 3.385 ;
        RECT  4.710 2.970 5.975 3.200 ;
        RECT  5.745 2.970 5.975 3.845 ;
        RECT  4.710 2.970 4.940 3.650 ;
        RECT  2.130 3.420 4.940 3.650 ;
        RECT  2.130 3.420 2.470 3.760 ;
        RECT  7.165 3.535 7.505 3.845 ;
        RECT  5.745 3.615 7.505 3.845 ;
        RECT  2.255 0.630 4.625 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  4.395 0.630 4.625 1.170 ;
        RECT  5.750 0.740 7.465 0.970 ;
        RECT  4.395 0.940 5.980 1.170 ;
        RECT  7.235 0.740 7.465 1.600 ;
        RECT  7.235 1.260 7.575 1.600 ;
        RECT  8.350 2.020 8.625 2.965 ;
        RECT  9.735 1.240 10.020 3.120 ;
        RECT  6.785 1.770 7.070 2.700 ;
        RECT  8.350 2.625 10.020 2.965 ;
        RECT  6.975 2.470 7.205 3.305 ;
        RECT  9.665 2.890 11.020 3.120 ;
        RECT  10.680 2.890 11.020 3.230 ;
        RECT  8.350 2.020 8.580 3.305 ;
        RECT  6.975 3.075 8.580 3.305 ;
        RECT  9.275 0.780 10.540 1.010 ;
        RECT  7.890 0.630 8.245 1.410 ;
        RECT  9.275 0.780 9.505 1.410 ;
        RECT  7.890 1.180 9.505 1.410 ;
        RECT  7.890 0.630 8.120 2.235 ;
        RECT  7.400 1.950 8.005 2.290 ;
        RECT  10.310 2.220 10.825 2.450 ;
        RECT  10.310 0.780 10.540 2.450 ;
        RECT  10.485 2.330 11.640 2.560 ;
        RECT  7.665 1.950 8.005 2.845 ;
        RECT  11.355 2.330 11.640 3.450 ;
        RECT  13.510 0.670 13.850 1.010 ;
        RECT  11.525 1.060 11.865 1.485 ;
        RECT  13.510 0.670 13.740 1.485 ;
        RECT  11.525 1.255 13.740 1.485 ;
        RECT  11.870 1.255 12.100 3.970 ;
        RECT  10.960 3.680 12.100 3.970 ;
        RECT  14.030 1.640 14.370 2.640 ;
        RECT  14.030 2.300 14.780 2.640 ;
        RECT  12.330 2.645 12.670 3.160 ;
        RECT  14.030 1.640 14.260 3.160 ;
        RECT  12.330 2.930 14.260 3.160 ;
        RECT  13.025 2.930 13.365 3.970 ;
        RECT  1.255 1.585 2.90 1.815 ;
        RECT  2.130 3.420 3.70 3.650 ;
        RECT  2.255 0.630 3.60 0.860 ;
        RECT  11.525 1.255 12.70 1.485 ;
    END
END SDFRSX1

MACRO SDFRSX0
    CLASS CORE ;
    FOREIGN SDFRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.489  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.480 2.640 14.995 3.240 ;
        RECT  14.670 1.170 14.995 3.240 ;
        RECT  14.560 1.170 14.995 1.510 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.628  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 1.640 14.365 2.020 ;
        RECT  13.615 2.620 14.215 2.960 ;
        RECT  13.985 0.630 14.215 2.960 ;
        RECT  13.305 0.630 14.215 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.315 2.415 2.545 ;
        RECT  0.705 2.255 1.045 2.545 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 2.225 8.850 2.675 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 2.250 12.690 2.660 ;
        END
    END SN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.480 3.470 14.820 5.280 ;
        RECT  13.160 4.165 13.500 5.280 ;
        RECT  11.735 3.630 12.020 5.280 ;
        RECT  8.960 3.630 9.300 5.280 ;
        RECT  8.025 3.880 8.365 5.280 ;
        RECT  4.830 3.910 5.115 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  14.560 -0.400 14.900 0.710 ;
        RECT  12.195 -0.400 12.535 0.930 ;
        RECT  10.110 -0.400 10.395 0.710 ;
        RECT  10.090 -0.400 10.395 0.675 ;
        RECT  8.165 -0.400 8.500 1.030 ;
        RECT  4.495 -0.400 4.835 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.555 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.815 ;
        RECT  2.930 1.585 3.270 1.960 ;
        RECT  0.245 1.795 1.320 2.025 ;
        RECT  0.245 1.795 0.475 3.380 ;
        RECT  0.245 2.885 1.305 3.215 ;
        RECT  0.245 2.885 0.785 3.380 ;
        RECT  3.505 1.805 5.295 2.035 ;
        RECT  3.505 1.805 3.970 2.095 ;
        RECT  5.010 1.805 5.295 2.205 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.525 1.230 6.430 1.540 ;
        RECT  3.965 2.325 4.250 2.665 ;
        RECT  3.965 2.435 5.755 2.665 ;
        RECT  5.525 1.230 5.755 3.220 ;
        RECT  5.520 2.435 5.755 3.220 ;
        RECT  5.520 2.990 6.235 3.220 ;
        RECT  6.005 2.990 6.235 3.790 ;
        RECT  6.005 3.450 6.345 3.790 ;
        RECT  4.370 3.450 5.575 3.680 ;
        RECT  4.370 3.450 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.345 3.450 5.575 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.765 3.880 7.105 4.250 ;
        RECT  5.345 4.020 7.105 4.250 ;
        RECT  5.065 0.770 7.255 1.000 ;
        RECT  1.980 0.980 2.320 1.355 ;
        RECT  5.065 0.770 5.295 1.355 ;
        RECT  1.980 1.125 5.295 1.355 ;
        RECT  6.915 0.770 7.255 1.570 ;
        RECT  5.985 2.440 6.325 2.760 ;
        RECT  7.675 2.330 8.025 2.695 ;
        RECT  5.985 2.530 6.805 2.760 ;
        RECT  9.190 1.230 9.420 3.190 ;
        RECT  9.190 2.850 10.250 3.190 ;
        RECT  7.795 2.905 10.250 3.190 ;
        RECT  6.575 2.530 6.805 3.650 ;
        RECT  7.795 2.330 8.025 3.650 ;
        RECT  6.575 3.420 8.025 3.650 ;
        RECT  8.730 0.770 9.880 1.000 ;
        RECT  8.730 0.770 8.960 1.590 ;
        RECT  7.615 1.360 8.960 1.590 ;
        RECT  5.985 1.770 6.270 2.110 ;
        RECT  7.615 1.360 7.955 2.030 ;
        RECT  5.985 1.800 7.955 2.030 ;
        RECT  9.650 0.770 9.880 2.290 ;
        RECT  5.985 1.800 7.445 2.110 ;
        RECT  9.650 2.060 10.265 2.290 ;
        RECT  9.925 2.170 10.935 2.400 ;
        RECT  7.215 1.800 7.445 3.190 ;
        RECT  7.215 2.880 7.535 3.190 ;
        RECT  10.705 2.170 10.935 3.440 ;
        RECT  7.215 2.905 7.565 3.190 ;
        RECT  10.705 3.100 11.045 3.440 ;
        RECT  10.965 1.110 11.505 1.450 ;
        RECT  12.590 3.060 12.910 3.400 ;
        RECT  11.275 3.170 12.910 3.400 ;
        RECT  11.275 1.110 11.505 3.970 ;
        RECT  10.255 3.670 11.505 3.970 ;
        RECT  13.305 1.310 13.645 2.320 ;
        RECT  11.925 1.670 13.645 2.020 ;
        RECT  13.140 1.980 13.755 2.320 ;
        RECT  13.140 1.670 13.370 3.900 ;
        RECT  12.360 3.650 13.370 3.900 ;
        RECT  12.360 3.650 12.745 3.970 ;
        RECT  0.980 1.585 2.60 1.815 ;
        RECT  1.995 3.710 3.80 3.940 ;
        RECT  5.065 0.770 6.30 1.000 ;
        RECT  1.980 1.125 4.40 1.355 ;
        RECT  7.795 2.905 9.60 3.190 ;
    END
END SDFRSX0

MACRO SDFRSQX4
    CLASS CORE ;
    FOREIGN SDFRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.075 2.250 17.415 4.100 ;
        RECT  15.635 2.250 17.415 2.630 ;
        RECT  16.560 1.230 16.900 2.630 ;
        RECT  15.635 2.250 15.975 4.100 ;
        RECT  15.540 0.700 15.770 2.480 ;
        RECT  15.240 0.700 15.770 1.040 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.760 1.640 14.365 2.020 ;
        RECT  13.760 1.640 14.105 2.200 ;
        END
    END SN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 1.660 9.500 2.100 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  17.120 -0.400 17.460 0.710 ;
        RECT  16.000 -0.400 16.340 0.710 ;
        RECT  13.190 -0.400 14.000 0.800 ;
        RECT  10.715 -0.400 11.000 1.370 ;
        RECT  8.820 -0.400 9.105 0.970 ;
        RECT  3.400 -0.400 5.150 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.355 2.860 16.695 5.280 ;
        RECT  14.875 4.140 15.215 5.280 ;
        RECT  13.590 2.890 13.930 5.280 ;
        RECT  11.370 3.965 11.710 5.280 ;
        RECT  8.975 2.910 9.260 5.280 ;
        RECT  4.795 3.965 5.135 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.585 5.740 1.875 ;
        RECT  5.400 1.585 5.740 2.265 ;
        RECT  3.895 1.585 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.025 1.190 6.800 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  6.025 1.190 6.255 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  6.025 2.935 6.450 3.275 ;
        RECT  4.630 3.045 6.450 3.275 ;
        RECT  6.830 2.980 7.170 3.735 ;
        RECT  2.020 3.505 7.170 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.380 0.730 7.260 0.960 ;
        RECT  2.255 0.940 5.610 1.170 ;
        RECT  7.030 0.730 7.260 1.660 ;
        RECT  7.030 1.320 7.615 1.660 ;
        RECT  9.335 0.775 10.485 1.005 ;
        RECT  7.490 0.735 8.360 1.090 ;
        RECT  8.000 0.735 8.360 1.430 ;
        RECT  9.335 0.775 9.565 1.430 ;
        RECT  8.000 1.200 9.565 1.430 ;
        RECT  10.255 0.775 10.485 1.960 ;
        RECT  10.255 1.730 11.910 1.960 ;
        RECT  11.570 1.730 11.910 2.070 ;
        RECT  8.000 0.735 8.285 2.940 ;
        RECT  6.485 1.840 6.795 2.195 ;
        RECT  6.485 1.965 7.770 2.195 ;
        RECT  9.795 1.240 10.025 2.680 ;
        RECT  9.795 2.340 10.740 2.680 ;
        RECT  12.240 1.540 12.525 2.680 ;
        RECT  8.515 2.450 12.525 2.680 ;
        RECT  9.640 2.450 9.980 2.860 ;
        RECT  7.430 1.965 7.770 3.400 ;
        RECT  8.515 2.450 8.745 3.400 ;
        RECT  7.430 3.170 8.745 3.400 ;
        RECT  9.640 2.450 9.870 3.855 ;
        RECT  10.840 3.505 12.180 3.735 ;
        RECT  11.950 3.505 12.180 4.100 ;
        RECT  9.640 3.625 11.070 3.855 ;
        RECT  11.950 3.760 12.460 4.100 ;
        RECT  11.810 0.970 12.150 1.310 ;
        RECT  11.810 1.080 12.985 1.310 ;
        RECT  14.505 2.320 14.845 2.660 ;
        RECT  12.755 2.430 14.845 2.660 ;
        RECT  12.755 1.080 12.985 3.220 ;
        RECT  10.180 2.990 12.985 3.220 ;
        RECT  12.360 2.990 12.700 3.330 ;
        RECT  10.180 2.990 10.520 3.395 ;
        RECT  13.215 1.180 15.010 1.410 ;
        RECT  14.670 1.180 15.010 1.700 ;
        RECT  13.215 1.180 13.500 1.530 ;
        RECT  14.670 1.470 15.310 1.700 ;
        RECT  15.080 1.470 15.310 3.120 ;
        RECT  14.315 2.890 15.310 3.120 ;
        RECT  14.315 2.890 14.655 3.730 ;
        RECT  1.145 1.585 2.70 1.815 ;
        RECT  2.020 3.505 6.60 3.735 ;
        RECT  2.255 0.940 4.60 1.170 ;
        RECT  8.515 2.450 11.90 2.680 ;
        RECT  12.755 2.430 13.70 2.660 ;
        RECT  10.180 2.990 11.00 3.220 ;
    END
END SDFRSQX4

MACRO SDFRSQX2
    CLASS CORE ;
    FOREIGN SDFRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.670 1.250 15.010 2.630 ;
        RECT  14.450 2.250 14.790 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.720 1.005 2.200 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 2.020 8.760 2.630 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.585 2.050 13.105 2.630 ;
        END
    END SN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.230 -0.400 15.570 0.720 ;
        RECT  14.110 -0.400 14.450 0.720 ;
        RECT  12.300 -0.400 12.645 1.090 ;
        RECT  9.910 -0.400 10.195 1.330 ;
        RECT  7.990 -0.400 8.275 1.330 ;
        RECT  4.530 -0.400 4.870 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.210 3.270 15.550 5.280 ;
        RECT  13.690 4.170 14.030 5.280 ;
        RECT  12.410 3.385 12.750 5.280 ;
        RECT  11.710 3.320 12.050 5.280 ;
        RECT  9.330 3.480 9.670 5.280 ;
        RECT  8.030 3.515 8.370 5.280 ;
        RECT  4.715 3.900 5.055 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.330 2.015 ;
        RECT  4.990 1.785 5.330 2.470 ;
        RECT  3.480 1.400 3.710 3.270 ;
        RECT  3.480 2.930 4.250 3.265 ;
        RECT  3.480 2.930 4.240 3.270 ;
        RECT  5.580 1.190 6.100 1.530 ;
        RECT  3.940 2.245 4.715 2.585 ;
        RECT  4.485 2.245 4.715 2.930 ;
        RECT  5.580 1.190 5.810 3.210 ;
        RECT  4.485 2.700 5.810 2.930 ;
        RECT  5.580 2.870 6.285 3.210 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  5.120 0.730 6.900 0.960 ;
        RECT  1.770 0.940 5.350 1.170 ;
        RECT  6.560 0.730 6.900 1.595 ;
        RECT  4.400 3.440 5.525 3.670 ;
        RECT  2.120 3.500 4.560 3.730 ;
        RECT  5.295 3.515 7.045 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  7.215 0.630 7.555 0.965 ;
        RECT  8.505 0.800 9.680 1.030 ;
        RECT  7.325 0.630 7.555 2.825 ;
        RECT  9.450 0.800 9.680 1.790 ;
        RECT  8.505 0.800 8.735 1.790 ;
        RECT  7.325 1.560 8.735 1.790 ;
        RECT  9.450 1.560 11.105 1.790 ;
        RECT  10.765 1.560 11.105 1.895 ;
        RECT  7.065 1.825 7.610 2.165 ;
        RECT  7.325 1.560 7.610 2.825 ;
        RECT  7.270 1.825 7.610 2.825 ;
        RECT  8.965 1.260 9.220 1.600 ;
        RECT  6.040 1.760 6.380 2.110 ;
        RECT  6.040 1.880 6.780 2.110 ;
        RECT  10.040 2.120 10.380 2.460 ;
        RECT  10.040 2.225 11.425 2.460 ;
        RECT  8.990 2.230 11.425 2.460 ;
        RECT  11.140 2.225 11.425 2.565 ;
        RECT  6.550 1.880 6.780 3.285 ;
        RECT  8.830 2.850 9.220 3.145 ;
        RECT  7.840 2.860 9.220 3.145 ;
        RECT  8.990 1.260 9.220 3.145 ;
        RECT  7.840 2.020 8.085 3.285 ;
        RECT  6.550 3.055 8.085 3.285 ;
        RECT  11.035 1.035 11.810 1.330 ;
        RECT  11.580 1.035 11.810 2.055 ;
        RECT  11.655 1.835 11.885 3.090 ;
        RECT  13.415 2.750 13.755 3.090 ;
        RECT  10.480 2.860 13.755 3.090 ;
        RECT  10.480 2.860 10.820 3.615 ;
        RECT  13.335 0.630 13.675 1.660 ;
        RECT  12.040 1.320 13.675 1.660 ;
        RECT  12.040 1.430 14.215 1.660 ;
        RECT  13.985 1.430 14.215 3.720 ;
        RECT  13.130 3.380 14.215 3.720 ;
        RECT  1.770 0.940 4.30 1.170 ;
        RECT  2.120 3.500 3.20 3.730 ;
        RECT  8.990 2.230 10.70 2.460 ;
        RECT  10.480 2.860 12.70 3.090 ;
        RECT  12.040 1.430 13.60 1.660 ;
    END
END SDFRSQX2

MACRO SDFRSQX1
    CLASS CORE ;
    FOREIGN SDFRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.855 1.660 9.385 2.120 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.250 14.995 2.630 ;
        RECT  14.410 3.625 14.845 3.965 ;
        RECT  14.615 0.700 14.845 3.965 ;
        RECT  14.410 0.700 14.845 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.670 3.995 2.030 4.250 ;
        RECT  1.670 3.960 2.015 4.250 ;
        RECT  1.670 3.470 1.900 4.250 ;
        RECT  1.410 3.470 1.900 3.815 ;
        RECT  1.385 3.470 1.900 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.940 2.800 3.655 3.190 ;
        RECT  2.940 2.045 3.170 3.190 ;
        RECT  0.575 2.045 3.170 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.805 2.710 3.190 ;
        RECT  2.370 2.505 2.710 3.190 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.075 2.250 13.735 2.700 ;
        END
    END SN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.130 -0.400 15.470 1.060 ;
        RECT  12.755 -0.400 13.095 1.025 ;
        RECT  10.770 -0.400 11.110 1.005 ;
        RECT  8.705 -0.400 9.045 0.970 ;
        RECT  5.170 -0.400 5.510 0.710 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  2.825 1.090 3.825 1.320 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.130 3.330 15.470 5.280 ;
        RECT  13.825 4.170 14.165 5.280 ;
        RECT  12.330 3.630 12.645 5.280 ;
        RECT  9.765 3.480 10.105 5.280 ;
        RECT  8.465 3.535 8.805 5.280 ;
        RECT  5.170 3.430 5.510 5.280 ;
        RECT  3.470 4.170 3.810 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.690 1.815 ;
        RECT  3.350 1.555 3.690 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  4.080 1.570 4.420 2.090 ;
        RECT  3.920 1.860 5.830 2.090 ;
        RECT  5.490 1.860 5.830 2.280 ;
        RECT  3.920 1.860 4.150 3.190 ;
        RECT  3.920 2.850 4.480 3.190 ;
        RECT  6.325 1.200 6.740 1.540 ;
        RECT  4.390 2.320 4.995 2.605 ;
        RECT  4.780 2.510 6.555 2.740 ;
        RECT  6.325 1.200 6.555 3.385 ;
        RECT  6.325 3.045 6.745 3.385 ;
        RECT  4.710 2.970 5.975 3.200 ;
        RECT  5.745 2.970 5.975 3.845 ;
        RECT  4.710 2.970 4.940 3.650 ;
        RECT  2.130 3.420 4.940 3.650 ;
        RECT  2.130 3.420 2.470 3.760 ;
        RECT  7.165 3.535 7.505 3.845 ;
        RECT  5.745 3.615 7.505 3.845 ;
        RECT  2.255 0.630 4.625 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  4.395 0.630 4.625 1.170 ;
        RECT  5.750 0.740 7.465 0.970 ;
        RECT  4.395 0.940 5.980 1.170 ;
        RECT  7.235 0.740 7.465 1.600 ;
        RECT  7.235 1.260 7.575 1.600 ;
        RECT  8.350 2.020 8.625 2.965 ;
        RECT  9.735 1.240 10.020 3.120 ;
        RECT  6.785 1.770 7.070 2.700 ;
        RECT  8.350 2.625 10.020 2.965 ;
        RECT  6.975 2.470 7.205 3.305 ;
        RECT  9.665 2.890 11.020 3.120 ;
        RECT  10.680 2.890 11.020 3.230 ;
        RECT  8.350 2.020 8.580 3.305 ;
        RECT  6.975 3.075 8.580 3.305 ;
        RECT  9.275 0.780 10.540 1.010 ;
        RECT  7.890 0.630 8.245 1.430 ;
        RECT  9.275 0.780 9.505 1.430 ;
        RECT  7.890 1.200 9.505 1.430 ;
        RECT  7.890 0.630 8.120 2.235 ;
        RECT  7.400 1.950 8.005 2.290 ;
        RECT  10.310 2.220 10.825 2.450 ;
        RECT  10.310 0.780 10.540 2.450 ;
        RECT  10.485 2.330 11.640 2.560 ;
        RECT  7.665 1.950 8.005 2.845 ;
        RECT  11.355 2.330 11.640 3.450 ;
        RECT  13.510 0.910 13.850 1.250 ;
        RECT  13.510 0.910 13.740 1.485 ;
        RECT  11.525 1.255 13.740 1.485 ;
        RECT  11.525 1.255 12.100 1.610 ;
        RECT  11.870 1.255 12.100 3.970 ;
        RECT  10.960 3.680 12.100 3.970 ;
        RECT  14.030 1.640 14.370 1.980 ;
        RECT  12.330 2.645 12.670 3.160 ;
        RECT  14.030 1.640 14.260 3.160 ;
        RECT  12.330 2.930 14.260 3.160 ;
        RECT  13.025 2.930 13.365 3.970 ;
        RECT  1.255 1.585 2.50 1.815 ;
        RECT  2.130 3.420 3.80 3.650 ;
        RECT  2.255 0.630 3.20 0.860 ;
        RECT  11.525 1.255 12.30 1.485 ;
    END
END SDFRSQX1

MACRO SDFRSQX0
    CLASS CORE ;
    FOREIGN SDFRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.560  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.340 2.250 13.745 3.050 ;
        RECT  13.515 0.630 13.745 3.050 ;
        RECT  12.990 0.630 13.745 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.555 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.255 2.120 8.700 2.670 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.980 2.240 12.585 2.705 ;
        END
    END SN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.950 4.020 13.290 5.280 ;
        RECT  11.395 3.910 11.680 5.280 ;
        RECT  8.760 3.630 9.100 5.280 ;
        RECT  8.025 3.880 8.365 5.280 ;
        RECT  4.830 3.910 5.115 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  11.880 -0.400 12.220 0.715 ;
        RECT  9.850 -0.400 10.190 0.710 ;
        RECT  7.900 -0.400 8.185 0.970 ;
        RECT  4.495 -0.400 4.835 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.235 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.505 1.805 5.295 2.095 ;
        RECT  5.010 1.805 5.295 2.205 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.525 1.230 6.430 1.540 ;
        RECT  3.965 2.325 4.250 2.665 ;
        RECT  3.965 2.435 5.755 2.665 ;
        RECT  5.525 1.230 5.755 3.220 ;
        RECT  5.520 2.435 5.755 3.220 ;
        RECT  5.520 2.990 6.235 3.220 ;
        RECT  6.005 2.990 6.235 3.790 ;
        RECT  6.005 3.450 6.345 3.790 ;
        RECT  4.370 3.450 5.575 3.680 ;
        RECT  4.370 3.450 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.345 3.450 5.575 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.765 3.880 7.105 4.250 ;
        RECT  5.345 4.020 7.105 4.250 ;
        RECT  5.065 0.630 7.110 0.860 ;
        RECT  6.770 0.630 7.110 0.970 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  5.065 0.630 5.295 1.355 ;
        RECT  1.980 1.125 5.295 1.355 ;
        RECT  8.875 1.230 9.160 1.570 ;
        RECT  5.985 2.440 6.325 2.760 ;
        RECT  7.675 2.355 8.025 2.695 ;
        RECT  5.985 2.530 6.805 2.760 ;
        RECT  8.930 2.710 10.050 2.940 ;
        RECT  9.710 2.600 10.050 2.940 ;
        RECT  8.930 1.230 9.160 3.190 ;
        RECT  7.795 2.905 9.160 3.190 ;
        RECT  6.575 2.530 6.805 3.650 ;
        RECT  7.795 2.355 8.025 3.650 ;
        RECT  6.575 3.420 8.025 3.650 ;
        RECT  8.415 0.770 9.620 1.000 ;
        RECT  8.415 0.770 8.645 1.490 ;
        RECT  7.390 1.250 8.645 1.490 ;
        RECT  9.390 0.770 9.620 2.160 ;
        RECT  7.390 1.250 7.730 2.030 ;
        RECT  5.985 1.770 7.445 2.110 ;
        RECT  9.390 1.930 10.130 2.160 ;
        RECT  9.790 2.040 10.595 2.270 ;
        RECT  7.215 1.770 7.445 3.190 ;
        RECT  7.215 2.880 7.535 3.190 ;
        RECT  10.365 2.040 10.595 3.415 ;
        RECT  7.215 2.905 7.565 3.190 ;
        RECT  10.365 3.075 10.705 3.415 ;
        RECT  10.650 1.110 11.165 1.450 ;
        RECT  10.935 2.990 12.630 3.330 ;
        RECT  10.935 1.110 11.165 3.970 ;
        RECT  9.990 3.645 11.165 3.970 ;
        RECT  12.990 1.310 13.285 1.900 ;
        RECT  11.395 1.670 13.090 2.010 ;
        RECT  11.395 1.670 11.705 2.310 ;
        RECT  12.860 1.670 13.090 3.790 ;
        RECT  12.140 3.560 13.090 3.790 ;
        RECT  12.140 3.560 12.480 3.880 ;
        RECT  0.980 1.585 2.20 1.960 ;
        RECT  1.995 3.710 3.50 3.940 ;
        RECT  5.065 0.630 6.10 0.860 ;
        RECT  1.980 1.125 4.40 1.355 ;
    END
END SDFRSQX0

MACRO SDFRRX4
    CLASS CORE ;
    FOREIGN SDFRRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.050 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  21.530 1.130 21.870 4.005 ;
        RECT  20.090 2.250 21.870 2.630 ;
        RECT  20.090 1.130 20.430 4.005 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.119  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.355 3.010 19.730 3.240 ;
        RECT  19.500 1.700 19.730 3.240 ;
        RECT  17.210 1.700 19.730 1.930 ;
        RECT  18.795 3.010 19.135 3.350 ;
        RECT  18.650 1.130 18.990 1.930 ;
        RECT  17.355 2.860 18.145 3.240 ;
        RECT  17.355 2.860 17.695 4.130 ;
        RECT  17.210 1.130 17.550 1.930 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.020 1.640 15.650 2.175 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.660 10.630 2.135 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 22.050 0.400 ;
        RECT  20.810 -0.400 21.150 1.470 ;
        RECT  19.370 -0.400 19.710 1.470 ;
        RECT  17.930 -0.400 18.270 1.470 ;
        RECT  15.670 -0.400 16.010 0.950 ;
        RECT  9.920 -0.400 10.205 0.970 ;
        RECT  4.775 -0.400 5.915 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 22.050 5.280 ;
        RECT  20.810 2.860 21.150 5.280 ;
        RECT  19.370 3.665 19.710 5.280 ;
        RECT  18.075 3.470 18.415 5.280 ;
        RECT  16.595 4.170 16.935 5.280 ;
        RECT  14.155 3.640 15.615 5.280 ;
        RECT  12.095 3.980 12.435 5.280 ;
        RECT  9.540 2.950 9.825 5.280 ;
        RECT  4.660 4.115 5.700 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 5.885 2.095 ;
        RECT  5.655 1.860 5.885 2.800 ;
        RECT  5.655 2.460 5.995 2.800 ;
        RECT  3.895 1.815 4.125 3.425 ;
        RECT  3.895 3.085 4.260 3.425 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 6.625 1.585 ;
        RECT  5.015 1.355 6.625 1.630 ;
        RECT  6.335 1.355 6.625 1.695 ;
        RECT  2.020 3.655 6.390 3.885 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  6.160 3.850 7.710 4.080 ;
        RECT  7.370 3.850 7.710 4.190 ;
        RECT  6.855 1.160 7.900 1.500 ;
        RECT  4.355 2.325 4.640 2.665 ;
        RECT  4.355 2.435 4.890 2.665 ;
        RECT  4.660 2.435 4.890 3.425 ;
        RECT  4.660 3.085 5.000 3.425 ;
        RECT  4.660 3.195 7.085 3.425 ;
        RECT  6.855 1.160 7.085 3.540 ;
        RECT  6.745 3.195 7.085 3.540 ;
        RECT  6.210 0.630 8.360 0.860 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.210 0.630 6.440 1.125 ;
        RECT  4.315 0.895 6.440 1.125 ;
        RECT  8.130 0.630 8.360 1.660 ;
        RECT  8.130 1.320 8.715 1.660 ;
        RECT  10.435 0.775 11.585 1.005 ;
        RECT  8.590 0.735 9.460 1.090 ;
        RECT  10.435 0.775 10.665 1.430 ;
        RECT  9.230 1.200 10.665 1.430 ;
        RECT  11.355 0.775 11.585 2.090 ;
        RECT  11.355 1.860 13.020 2.090 ;
        RECT  9.230 0.735 9.460 2.150 ;
        RECT  8.620 1.920 9.460 2.150 ;
        RECT  12.680 1.860 13.020 2.200 ;
        RECT  8.620 1.920 8.850 3.580 ;
        RECT  8.510 3.235 8.850 3.580 ;
        RECT  13.350 1.670 13.690 2.010 ;
        RECT  7.315 1.800 7.625 2.160 ;
        RECT  10.895 1.240 11.125 2.680 ;
        RECT  10.895 2.340 11.485 2.680 ;
        RECT  13.350 1.670 13.580 2.680 ;
        RECT  9.080 2.450 13.580 2.680 ;
        RECT  7.395 1.800 7.625 3.205 ;
        RECT  7.395 2.865 8.280 3.205 ;
        RECT  10.205 2.450 10.545 3.915 ;
        RECT  11.565 3.520 12.895 3.750 ;
        RECT  12.665 3.520 12.895 4.180 ;
        RECT  10.205 3.685 11.795 3.915 ;
        RECT  8.050 2.865 8.280 4.185 ;
        RECT  12.665 3.840 13.185 4.180 ;
        RECT  9.080 2.450 9.310 4.185 ;
        RECT  8.050 3.955 9.310 4.185 ;
        RECT  11.815 0.630 15.210 0.860 ;
        RECT  14.385 0.630 15.210 0.950 ;
        RECT  11.815 0.630 12.110 1.500 ;
        RECT  12.920 1.090 14.150 1.375 ;
        RECT  15.950 2.370 16.290 2.710 ;
        RECT  13.920 2.480 16.290 2.710 ;
        RECT  14.715 2.480 15.055 3.050 ;
        RECT  13.920 1.090 14.150 3.215 ;
        RECT  10.905 2.985 14.150 3.215 ;
        RECT  10.905 2.985 11.245 3.455 ;
        RECT  13.125 2.985 13.465 3.610 ;
        RECT  16.430 1.070 16.770 1.410 ;
        RECT  14.380 1.180 16.770 1.410 ;
        RECT  14.380 1.180 14.720 1.675 ;
        RECT  16.540 2.310 19.270 2.540 ;
        RECT  18.985 2.310 19.270 2.650 ;
        RECT  16.540 1.070 16.770 3.170 ;
        RECT  16.035 2.940 16.770 3.170 ;
        RECT  16.035 2.940 16.375 3.760 ;
        RECT  1.145 1.585 2.80 1.815 ;
        RECT  1.605 1.125 3.40 1.355 ;
        RECT  3.855 1.355 5.40 1.585 ;
        RECT  2.020 3.655 5.30 3.885 ;
        RECT  4.660 3.195 6.20 3.425 ;
        RECT  6.210 0.630 7.50 0.860 ;
        RECT  2.255 0.630 3.00 0.895 ;
        RECT  4.315 0.895 5.40 1.125 ;
        RECT  9.080 2.450 12.80 2.680 ;
        RECT  11.815 0.630 14.40 0.860 ;
        RECT  13.920 2.480 15.90 2.710 ;
        RECT  10.905 2.985 13.40 3.215 ;
        RECT  14.380 1.180 15.90 1.410 ;
        RECT  16.540 2.310 18.30 2.540 ;
    END
END SDFRRX4

MACRO SDFRRX2
    CLASS CORE ;
    FOREIGN SDFRRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.270 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.020 0.820 16.255 3.240 ;
        RECT  15.710 2.860 16.105 3.830 ;
        RECT  15.870 0.820 16.255 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.250 9.700 2.630 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.200 2.110 13.735 2.675 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.135 1.230 17.530 2.020 ;
        RECT  17.030 2.640 17.370 3.550 ;
        RECT  17.135 1.230 17.370 3.550 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.270 0.400 ;
        RECT  17.750 -0.400 18.090 0.710 ;
        RECT  16.630 -0.400 16.970 0.710 ;
        RECT  15.110 -0.400 15.450 0.970 ;
        RECT  14.005 -0.400 14.345 1.220 ;
        RECT  9.035 -0.400 9.320 1.330 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.270 5.280 ;
        RECT  17.750 2.640 18.090 5.280 ;
        RECT  16.470 3.950 16.810 5.280 ;
        RECT  14.950 3.775 15.290 5.280 ;
        RECT  12.745 3.365 13.085 5.280 ;
        RECT  9.895 3.525 10.235 5.280 ;
        RECT  8.595 3.810 8.935 5.280 ;
        RECT  4.655 3.960 5.645 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.685 ;
        RECT  4.710 1.400 5.915 1.685 ;
        RECT  4.135 1.550 4.475 2.180 ;
        RECT  3.895 1.950 6.165 2.180 ;
        RECT  5.825 1.950 6.165 2.375 ;
        RECT  3.895 1.950 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.805 1.260 7.145 1.600 ;
        RECT  6.495 1.370 7.145 1.600 ;
        RECT  4.415 2.410 5.045 2.750 ;
        RECT  4.705 2.410 5.045 3.270 ;
        RECT  6.495 1.370 6.725 3.270 ;
        RECT  4.705 3.040 6.875 3.270 ;
        RECT  6.535 3.040 6.875 3.625 ;
        RECT  2.120 3.500 6.305 3.730 ;
        RECT  6.075 3.500 6.305 4.125 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  7.295 3.810 7.635 4.125 ;
        RECT  6.075 3.895 7.635 4.125 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.800 7.945 1.030 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  7.605 0.800 7.945 1.600 ;
        RECT  9.550 0.800 10.700 1.030 ;
        RECT  8.260 0.630 8.600 1.790 ;
        RECT  10.470 0.800 10.700 1.790 ;
        RECT  9.550 0.800 9.780 1.790 ;
        RECT  8.260 1.560 9.780 1.790 ;
        RECT  10.470 1.560 12.125 1.790 ;
        RECT  11.785 1.560 12.125 1.895 ;
        RECT  8.260 0.630 8.490 2.060 ;
        RECT  7.755 1.830 8.490 2.060 ;
        RECT  7.755 1.830 8.165 2.170 ;
        RECT  7.825 1.830 8.165 3.120 ;
        RECT  6.955 1.910 7.335 2.220 ;
        RECT  10.810 2.225 11.150 2.565 ;
        RECT  10.810 2.330 12.320 2.565 ;
        RECT  11.995 2.225 12.320 2.565 ;
        RECT  10.010 2.335 12.320 2.565 ;
        RECT  8.425 2.305 8.715 3.165 ;
        RECT  10.010 1.260 10.240 3.165 ;
        RECT  8.425 2.860 10.240 3.165 ;
        RECT  7.105 1.910 7.335 3.580 ;
        RECT  8.425 2.305 8.670 3.580 ;
        RECT  7.105 3.350 8.670 3.580 ;
        RECT  10.930 0.630 13.625 0.860 ;
        RECT  13.285 0.630 13.625 1.105 ;
        RECT  10.930 0.630 11.215 1.330 ;
        RECT  12.055 1.090 12.780 1.330 ;
        RECT  13.965 2.400 14.935 2.740 ;
        RECT  12.550 1.090 12.780 3.135 ;
        RECT  13.965 2.400 14.195 3.135 ;
        RECT  11.300 2.905 14.195 3.135 ;
        RECT  11.300 2.905 11.640 3.690 ;
        RECT  13.465 2.905 13.805 4.175 ;
        RECT  13.010 1.380 13.355 1.720 ;
        RECT  13.010 1.490 15.145 1.720 ;
        RECT  14.805 1.490 15.145 2.100 ;
        RECT  14.805 1.870 15.665 2.100 ;
        RECT  15.165 1.870 15.665 2.210 ;
        RECT  15.165 1.870 15.395 3.310 ;
        RECT  14.425 2.970 15.395 3.310 ;
        RECT  1.255 1.585 2.20 1.815 ;
        RECT  2.825 1.090 3.80 1.320 ;
        RECT  1.715 1.125 2.60 1.355 ;
        RECT  3.895 1.950 5.30 2.180 ;
        RECT  4.705 3.040 5.20 3.270 ;
        RECT  2.120 3.500 5.50 3.730 ;
        RECT  2.255 0.630 4.00 0.860 ;
        RECT  10.010 2.335 11.40 2.565 ;
        RECT  10.930 0.630 12.60 0.860 ;
        RECT  11.300 2.905 13.50 3.135 ;
        RECT  13.010 1.490 14.10 1.720 ;
    END
END SDFRRX2

MACRO SDFRRX1
    CLASS CORE ;
    FOREIGN SDFRRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.865 0.940 16.255 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.245 1.640 15.635 2.020 ;
        RECT  14.735 2.870 15.480 3.100 ;
        RECT  15.245 1.640 15.480 3.100 ;
        RECT  15.245 1.260 15.475 3.100 ;
        RECT  14.680 1.260 15.475 1.490 ;
        RECT  14.420 3.780 14.965 4.120 ;
        RECT  14.735 2.870 14.965 4.120 ;
        RECT  14.680 0.700 14.910 1.490 ;
        RECT  14.420 0.700 14.910 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.665 3.995 2.030 4.250 ;
        RECT  1.665 3.960 2.010 4.250 ;
        RECT  1.665 3.470 1.895 4.250 ;
        RECT  1.410 3.470 1.895 3.815 ;
        RECT  1.385 3.470 1.895 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.970 2.800 3.655 3.240 ;
        RECT  2.970 2.045 3.200 3.240 ;
        RECT  0.575 2.045 3.200 2.275 ;
        RECT  0.575 1.660 0.860 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.030 1.660 9.480 2.130 ;
        RECT  8.945 1.660 9.480 2.030 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.745 2.170 13.280 2.630 ;
        END
    END RN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.140 -0.400 15.480 1.030 ;
        RECT  13.460 -0.400 13.800 0.950 ;
        RECT  8.820 -0.400 9.105 0.970 ;
        RECT  4.815 -0.400 5.155 0.655 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.195 3.330 15.480 5.280 ;
        RECT  12.740 3.820 13.085 5.280 ;
        RECT  10.125 3.480 10.465 5.280 ;
        RECT  8.825 3.535 9.165 5.280 ;
        RECT  8.870 3.530 9.165 5.280 ;
        RECT  4.910 3.845 5.870 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.130 0.900 1.430 ;
        RECT  0.115 1.200 1.485 1.430 ;
        RECT  1.255 1.200 1.485 1.815 ;
        RECT  1.255 1.585 3.665 1.815 ;
        RECT  3.380 1.555 3.665 1.895 ;
        RECT  0.115 1.130 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.125 1.320 ;
        RECT  3.485 1.090 4.125 1.325 ;
        RECT  3.895 1.090 4.125 1.580 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  3.895 1.345 5.685 1.580 ;
        RECT  5.345 1.345 5.685 1.650 ;
        RECT  3.900 1.810 5.170 2.040 ;
        RECT  5.000 1.880 5.965 2.220 ;
        RECT  3.900 1.810 4.220 3.425 ;
        RECT  6.320 1.230 6.915 1.540 ;
        RECT  4.450 2.325 4.760 3.155 ;
        RECT  6.320 1.230 6.550 3.155 ;
        RECT  4.450 2.870 6.550 3.155 ;
        RECT  4.450 2.925 7.100 3.155 ;
        RECT  6.760 2.925 7.100 3.385 ;
        RECT  2.255 0.630 4.585 0.860 ;
        RECT  4.355 0.630 4.585 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.740 0.770 7.660 1.000 ;
        RECT  4.355 0.885 5.970 1.115 ;
        RECT  7.375 0.770 7.660 1.600 ;
        RECT  2.125 3.420 2.410 3.760 ;
        RECT  4.450 3.385 6.330 3.615 ;
        RECT  2.125 3.530 3.580 3.760 ;
        RECT  7.520 3.535 7.860 3.845 ;
        RECT  6.100 3.615 7.860 3.845 ;
        RECT  4.450 3.385 4.680 3.885 ;
        RECT  3.365 3.655 4.680 3.885 ;
        RECT  8.350 2.020 8.715 2.360 ;
        RECT  8.525 2.225 8.820 2.440 ;
        RECT  6.780 1.800 7.065 2.695 ;
        RECT  9.795 1.240 10.025 3.120 ;
        RECT  6.780 2.465 7.565 2.695 ;
        RECT  8.590 2.625 10.025 2.965 ;
        RECT  7.335 2.465 7.565 3.305 ;
        RECT  9.795 2.890 11.375 3.120 ;
        RECT  11.035 2.890 11.375 3.230 ;
        RECT  8.590 2.225 8.820 3.305 ;
        RECT  7.335 3.075 8.820 3.305 ;
        RECT  9.335 0.780 10.485 1.010 ;
        RECT  8.020 0.630 8.360 1.430 ;
        RECT  9.335 0.780 9.565 1.430 ;
        RECT  7.890 1.200 9.565 1.430 ;
        RECT  7.890 1.200 8.120 2.845 ;
        RECT  7.525 1.830 8.120 2.170 ;
        RECT  10.255 0.780 10.485 2.450 ;
        RECT  10.255 2.220 11.095 2.450 ;
        RECT  10.755 2.330 11.840 2.560 ;
        RECT  7.885 1.830 8.120 2.845 ;
        RECT  7.885 2.590 8.350 2.845 ;
        RECT  7.885 2.605 8.360 2.845 ;
        RECT  11.610 2.330 11.840 3.450 ;
        RECT  11.610 3.110 12.050 3.450 ;
        RECT  10.715 0.630 13.040 0.860 ;
        RECT  10.715 0.630 11.000 1.005 ;
        RECT  12.700 0.630 13.040 1.220 ;
        RECT  11.470 1.090 11.810 1.430 ;
        RECT  11.470 1.200 12.300 1.430 ;
        RECT  12.070 1.200 12.300 2.810 ;
        RECT  12.280 2.580 12.515 3.145 ;
        RECT  13.760 2.740 14.045 3.090 ;
        RECT  12.280 2.860 14.045 3.090 ;
        RECT  12.280 2.860 13.580 3.145 ;
        RECT  12.280 2.580 12.510 3.970 ;
        RECT  11.320 3.680 12.510 3.970 ;
        RECT  12.530 1.495 12.815 1.835 ;
        RECT  12.530 1.605 14.400 1.835 ;
        RECT  14.060 1.660 14.510 1.945 ;
        RECT  14.275 1.660 14.510 2.640 ;
        RECT  14.275 2.300 14.775 2.640 ;
        RECT  14.275 1.660 14.505 3.550 ;
        RECT  13.820 3.320 14.505 3.550 ;
        RECT  13.820 3.320 14.050 4.160 ;
        RECT  13.710 3.820 14.050 4.160 ;
        RECT  1.255 1.585 2.40 1.815 ;
        RECT  4.450 2.870 5.60 3.155 ;
        RECT  4.450 2.925 6.40 3.155 ;
        RECT  2.255 0.630 3.80 0.860 ;
        RECT  10.715 0.630 12.40 0.860 ;
    END
END SDFRRX1

MACRO SDFRRX0
    CLASS CORE ;
    FOREIGN SDFRRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.225 1.260 15.625 4.150 ;
        RECT  15.100 1.260 15.625 1.600 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.550  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.300 2.860 14.995 3.350 ;
        RECT  14.765 1.830 14.995 3.350 ;
        RECT  14.515 1.830 14.995 2.060 ;
        RECT  14.515 0.630 14.745 2.060 ;
        RECT  14.200 0.630 14.745 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.265 2.415 2.550 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.830 2.215 9.325 2.720 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.610 2.250 13.105 2.895 ;
        END
    END RN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  14.300 3.810 14.700 5.280 ;
        RECT  12.285 3.910 12.620 5.280 ;
        RECT  9.510 3.650 9.850 5.280 ;
        RECT  8.310 3.910 8.650 5.280 ;
        RECT  4.830 3.865 5.170 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.100 -0.400 15.440 0.800 ;
        RECT  13.400 -0.400 13.740 0.950 ;
        RECT  8.615 -0.400 8.900 1.400 ;
        RECT  4.485 -0.400 4.825 0.655 ;
        RECT  0.180 -0.400 0.520 1.575 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.815 ;
        RECT  2.930 1.585 3.270 1.960 ;
        RECT  0.245 1.805 1.320 2.035 ;
        RECT  0.245 1.805 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.230 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  3.500 1.345 5.425 1.575 ;
        RECT  3.505 1.805 5.520 2.090 ;
        RECT  5.235 1.805 5.520 2.160 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.750 1.230 6.655 1.540 ;
        RECT  3.965 2.325 4.950 2.665 ;
        RECT  4.605 2.325 4.950 3.175 ;
        RECT  4.605 2.945 5.980 3.175 ;
        RECT  5.750 1.230 5.980 3.175 ;
        RECT  5.780 3.060 6.500 3.290 ;
        RECT  6.270 3.060 6.500 3.790 ;
        RECT  6.270 3.450 6.610 3.790 ;
        RECT  4.370 3.455 5.605 3.635 ;
        RECT  4.370 3.405 5.580 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.420 3.485 5.650 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.030 3.910 7.370 4.250 ;
        RECT  5.420 4.020 7.370 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  3.960 0.630 4.190 1.115 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  5.290 0.770 7.455 1.000 ;
        RECT  3.960 0.885 5.520 1.115 ;
        RECT  7.115 0.770 7.455 1.570 ;
        RECT  6.210 2.490 6.545 2.830 ;
        RECT  7.875 2.360 8.310 2.700 ;
        RECT  6.210 2.530 7.075 2.830 ;
        RECT  8.910 2.990 9.250 3.395 ;
        RECT  9.590 1.230 9.820 3.395 ;
        RECT  10.460 3.055 10.800 3.395 ;
        RECT  8.080 3.165 10.800 3.395 ;
        RECT  6.845 2.530 7.075 3.680 ;
        RECT  8.080 2.360 8.310 3.680 ;
        RECT  6.845 3.450 8.310 3.680 ;
        RECT  9.130 0.770 10.280 1.000 ;
        RECT  7.815 1.230 8.155 1.870 ;
        RECT  7.815 1.640 9.360 1.870 ;
        RECT  9.130 0.770 9.360 1.870 ;
        RECT  6.210 1.820 8.045 2.110 ;
        RECT  6.210 1.820 7.645 2.160 ;
        RECT  10.050 0.770 10.280 2.425 ;
        RECT  10.050 2.195 10.800 2.425 ;
        RECT  10.460 2.305 11.485 2.535 ;
        RECT  7.415 1.820 7.645 3.220 ;
        RECT  7.415 2.925 7.825 3.220 ;
        RECT  11.255 2.305 11.485 3.460 ;
        RECT  7.415 2.930 7.850 3.220 ;
        RECT  11.255 3.120 11.595 3.460 ;
        RECT  10.510 0.635 12.860 0.865 ;
        RECT  10.510 0.635 10.850 0.975 ;
        RECT  12.520 0.635 12.860 0.975 ;
        RECT  11.485 1.175 12.055 1.515 ;
        RECT  11.825 3.125 13.610 3.465 ;
        RECT  10.805 3.660 11.140 3.990 ;
        RECT  10.805 3.675 11.145 3.990 ;
        RECT  11.825 1.175 12.055 3.990 ;
        RECT  10.805 3.705 12.055 3.990 ;
        RECT  13.840 1.410 14.285 1.750 ;
        RECT  12.450 1.735 14.070 2.020 ;
        RECT  13.840 2.290 14.535 2.630 ;
        RECT  13.840 1.410 14.070 4.175 ;
        RECT  13.195 3.835 14.070 4.175 ;
        RECT  0.980 1.585 2.40 1.815 ;
        RECT  1.445 1.125 2.30 1.355 ;
        RECT  3.505 1.805 4.20 2.090 ;
        RECT  1.995 3.710 3.80 3.940 ;
        RECT  1.980 0.630 3.80 0.860 ;
        RECT  5.290 0.770 6.80 1.000 ;
        RECT  8.080 3.165 9.30 3.395 ;
        RECT  10.510 0.635 11.70 0.865 ;
    END
END SDFRRX0

MACRO SDFRRSX4
    CLASS CORE ;
    FOREIGN SDFRRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.680 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.105  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  22.160 1.130 22.500 3.295 ;
        RECT  20.830 2.250 22.500 2.630 ;
        RECT  20.830 2.250 21.205 3.295 ;
        RECT  20.830 1.130 21.060 3.295 ;
        RECT  20.720 1.130 21.060 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.135  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.155 3.010 20.585 3.240 ;
        RECT  20.355 1.700 20.585 3.240 ;
        RECT  18.055 1.700 20.585 1.930 ;
        RECT  19.595 3.010 19.935 3.350 ;
        RECT  19.280 1.130 19.620 1.930 ;
        RECT  18.155 2.860 18.775 3.240 ;
        RECT  18.155 2.860 18.495 4.030 ;
        RECT  18.055 1.130 18.285 1.930 ;
        RECT  17.840 1.130 18.285 1.470 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.225 1.640 16.885 2.020 ;
        RECT  16.225 1.640 16.565 2.130 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.185 2.190 15.685 2.690 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 1.660 11.015 2.100 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 22.680 0.400 ;
        RECT  21.440 -0.400 21.780 1.470 ;
        RECT  20.000 -0.400 20.340 1.470 ;
        RECT  18.560 -0.400 18.900 1.470 ;
        RECT  15.945 -0.400 16.285 0.950 ;
        RECT  10.350 -0.400 10.635 0.970 ;
        RECT  4.775 -0.400 6.345 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 22.680 5.280 ;
        RECT  21.520 3.530 21.860 5.280 ;
        RECT  20.145 3.685 20.485 5.280 ;
        RECT  18.875 3.470 19.215 5.280 ;
        RECT  17.395 4.070 17.735 5.280 ;
        RECT  14.955 3.910 16.415 5.280 ;
        RECT  12.655 3.965 12.995 5.280 ;
        RECT  10.235 2.910 10.535 5.280 ;
        RECT  4.830 3.965 6.300 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 6.485 2.095 ;
        RECT  6.255 1.860 6.485 2.800 ;
        RECT  6.255 2.460 6.595 2.800 ;
        RECT  3.895 1.815 4.125 3.370 ;
        RECT  3.895 3.085 4.260 3.370 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 7.055 1.585 ;
        RECT  5.445 1.355 7.055 1.630 ;
        RECT  6.765 1.355 7.055 1.695 ;
        RECT  7.285 1.160 8.330 1.500 ;
        RECT  4.355 2.325 5.600 2.665 ;
        RECT  5.260 2.325 5.600 3.275 ;
        RECT  7.285 1.160 7.515 3.540 ;
        RECT  5.260 3.045 7.515 3.275 ;
        RECT  7.200 3.200 7.545 3.540 ;
        RECT  4.450 3.505 6.820 3.735 ;
        RECT  6.590 3.505 6.820 4.000 ;
        RECT  2.020 3.600 4.640 3.830 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  8.010 2.980 8.350 4.000 ;
        RECT  6.590 3.770 8.350 4.000 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.640 0.700 8.790 0.930 ;
        RECT  4.315 0.895 6.870 1.125 ;
        RECT  8.560 0.700 8.790 1.660 ;
        RECT  8.560 1.320 9.145 1.660 ;
        RECT  10.865 0.775 12.015 1.005 ;
        RECT  9.020 0.735 9.890 1.090 ;
        RECT  10.865 0.775 11.095 1.430 ;
        RECT  9.660 1.200 11.095 1.430 ;
        RECT  11.785 0.775 12.015 2.090 ;
        RECT  11.785 1.860 13.450 2.090 ;
        RECT  9.660 0.735 9.890 2.150 ;
        RECT  9.260 1.920 9.890 2.150 ;
        RECT  13.110 1.860 13.450 2.200 ;
        RECT  9.260 1.920 9.545 3.195 ;
        RECT  13.780 1.670 14.120 2.010 ;
        RECT  7.745 1.890 9.030 2.120 ;
        RECT  7.745 1.815 8.055 2.175 ;
        RECT  11.325 1.240 11.555 2.680 ;
        RECT  11.325 2.340 12.025 2.680 ;
        RECT  13.780 1.670 14.010 2.680 ;
        RECT  9.775 2.450 14.010 2.680 ;
        RECT  10.915 2.450 11.255 2.860 ;
        RECT  8.690 1.890 9.030 3.655 ;
        RECT  10.915 2.450 11.145 3.855 ;
        RECT  9.775 2.450 10.005 3.655 ;
        RECT  8.690 3.425 10.005 3.655 ;
        RECT  12.125 3.505 13.635 3.735 ;
        RECT  13.405 3.505 13.635 4.100 ;
        RECT  10.915 3.625 12.355 3.855 ;
        RECT  13.405 3.760 13.745 4.100 ;
        RECT  12.245 0.630 15.485 0.860 ;
        RECT  14.675 0.630 15.485 0.950 ;
        RECT  12.245 0.630 12.540 1.500 ;
        RECT  13.350 1.100 13.690 1.440 ;
        RECT  13.350 1.210 14.580 1.440 ;
        RECT  17.025 2.270 17.365 2.610 ;
        RECT  16.375 2.380 17.365 2.610 ;
        RECT  14.350 1.210 14.580 3.275 ;
        RECT  16.375 2.380 16.605 3.275 ;
        RECT  11.465 3.045 16.605 3.275 ;
        RECT  15.515 3.045 15.855 3.385 ;
        RECT  11.465 3.045 11.805 3.395 ;
        RECT  13.975 3.045 14.265 3.780 ;
        RECT  14.810 1.180 17.480 1.410 ;
        RECT  14.810 1.180 15.150 1.675 ;
        RECT  17.140 1.180 17.480 2.040 ;
        RECT  17.140 1.810 17.825 2.040 ;
        RECT  17.595 2.250 20.125 2.480 ;
        RECT  19.785 2.250 20.125 2.590 ;
        RECT  17.595 1.810 17.825 3.070 ;
        RECT  16.835 2.840 17.825 3.070 ;
        RECT  16.835 2.840 17.175 3.660 ;
        RECT  1.145 1.585 2.30 1.815 ;
        RECT  3.895 1.860 5.70 2.095 ;
        RECT  1.605 1.125 3.10 1.355 ;
        RECT  3.855 1.355 6.30 1.585 ;
        RECT  5.260 3.045 6.20 3.275 ;
        RECT  4.450 3.505 5.80 3.735 ;
        RECT  2.020 3.600 3.60 3.830 ;
        RECT  2.255 0.630 3.60 0.895 ;
        RECT  6.640 0.700 7.90 0.930 ;
        RECT  4.315 0.895 5.80 1.125 ;
        RECT  9.775 2.450 13.20 2.680 ;
        RECT  12.245 0.630 14.80 0.860 ;
        RECT  11.465 3.045 15.30 3.275 ;
        RECT  14.810 1.180 16.70 1.410 ;
        RECT  17.595 2.250 19.30 2.480 ;
    END
END SDFRRSX4

MACRO SDFRRSX2
    CLASS CORE ;
    FOREIGN SDFRRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.650 0.820 16.885 3.240 ;
        RECT  16.340 2.860 16.735 4.180 ;
        RECT  16.500 0.820 16.885 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.020 10.040 2.630 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 2.035 14.125 2.375 ;
        RECT  13.355 2.035 13.735 2.630 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.050 14.995 2.630 ;
        RECT  14.475 2.050 14.995 2.395 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.765 1.230 18.160 2.020 ;
        RECT  17.660 2.640 18.000 3.550 ;
        RECT  17.765 1.230 18.000 3.550 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  18.380 -0.400 18.720 0.710 ;
        RECT  17.260 -0.400 17.600 0.710 ;
        RECT  15.740 -0.400 16.080 0.970 ;
        RECT  14.395 -0.400 14.735 0.890 ;
        RECT  9.385 -0.400 9.670 1.330 ;
        RECT  5.630 -0.400 5.920 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  18.380 2.640 18.720 5.280 ;
        RECT  17.100 3.950 17.440 5.280 ;
        RECT  15.580 4.170 15.920 5.280 ;
        RECT  14.260 3.910 14.600 5.280 ;
        RECT  13.120 3.825 13.460 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.965 3.900 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.265 1.630 ;
        RECT  4.135 1.550 4.475 2.090 ;
        RECT  3.895 1.860 6.545 2.090 ;
        RECT  6.205 1.860 6.545 2.375 ;
        RECT  3.895 1.860 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.850 1.190 7.495 1.530 ;
        RECT  4.355 2.320 5.645 2.635 ;
        RECT  6.850 1.190 7.080 3.210 ;
        RECT  5.305 2.320 5.645 3.210 ;
        RECT  6.850 2.870 7.510 3.210 ;
        RECT  5.305 2.980 7.510 3.210 ;
        RECT  4.505 3.440 6.705 3.670 ;
        RECT  2.120 3.500 4.735 3.730 ;
        RECT  7.930 3.535 8.270 3.845 ;
        RECT  6.475 3.615 8.270 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.150 0.725 8.295 0.955 ;
        RECT  5.170 0.940 6.380 1.170 ;
        RECT  7.955 0.725 8.295 1.600 ;
        RECT  9.900 0.800 11.050 1.030 ;
        RECT  8.570 0.630 8.950 1.790 ;
        RECT  10.820 0.800 11.050 1.790 ;
        RECT  9.900 0.800 10.130 1.790 ;
        RECT  8.570 1.560 10.130 1.790 ;
        RECT  10.820 1.560 12.475 1.790 ;
        RECT  12.135 1.560 12.475 1.895 ;
        RECT  8.240 2.020 8.800 2.360 ;
        RECT  8.570 0.630 8.800 2.845 ;
        RECT  8.460 2.020 8.800 2.845 ;
        RECT  7.310 1.795 7.650 2.115 ;
        RECT  7.310 1.885 7.970 2.115 ;
        RECT  11.245 2.120 11.585 2.460 ;
        RECT  11.245 2.225 12.630 2.460 ;
        RECT  10.360 2.230 12.630 2.460 ;
        RECT  12.345 2.225 12.630 2.565 ;
        RECT  9.030 2.020 9.345 3.145 ;
        RECT  7.740 1.885 7.970 3.305 ;
        RECT  9.030 2.860 10.590 3.145 ;
        RECT  10.360 1.260 10.590 3.145 ;
        RECT  7.740 3.075 9.260 3.305 ;
        RECT  11.280 0.630 13.975 0.860 ;
        RECT  13.635 0.630 13.975 1.105 ;
        RECT  11.280 0.630 11.565 1.330 ;
        RECT  12.405 1.090 13.090 1.330 ;
        RECT  12.860 1.090 13.090 3.090 ;
        RECT  13.965 2.605 14.305 3.090 ;
        RECT  15.225 2.750 15.565 3.090 ;
        RECT  11.725 2.860 15.565 3.090 ;
        RECT  11.725 2.860 12.065 3.615 ;
        RECT  13.355 1.380 13.705 1.720 ;
        RECT  13.355 1.490 15.765 1.720 ;
        RECT  15.425 1.490 15.765 2.210 ;
        RECT  15.425 1.870 16.285 2.210 ;
        RECT  15.795 1.870 16.025 3.720 ;
        RECT  15.020 3.380 16.025 3.720 ;
        RECT  1.255 1.585 2.70 1.815 ;
        RECT  2.825 1.090 3.90 1.320 ;
        RECT  1.715 1.125 2.70 1.355 ;
        RECT  3.895 1.860 5.80 2.090 ;
        RECT  5.305 2.980 6.30 3.210 ;
        RECT  4.505 3.440 5.20 3.670 ;
        RECT  2.120 3.500 3.80 3.730 ;
        RECT  2.255 0.630 4.60 0.860 ;
        RECT  6.150 0.725 7.40 0.955 ;
        RECT  10.360 2.230 11.90 2.460 ;
        RECT  11.280 0.630 12.40 0.860 ;
        RECT  11.725 2.860 14.60 3.090 ;
        RECT  13.355 1.490 14.50 1.720 ;
    END
END SDFRRSX2

MACRO SDFRRSX1
    CLASS CORE ;
    FOREIGN SDFRRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 2.860 17.515 3.240 ;
        RECT  17.120 0.940 17.460 1.280 ;
        RECT  17.120 2.860 17.450 4.180 ;
        RECT  17.120 0.940 17.350 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.425 1.640 16.885 2.020 ;
        RECT  15.885 2.870 16.655 3.100 ;
        RECT  16.425 1.235 16.655 3.100 ;
        RECT  15.840 1.235 16.655 1.465 ;
        RECT  15.670 3.680 16.115 3.965 ;
        RECT  15.885 2.870 16.115 3.965 ;
        RECT  15.840 0.700 16.070 1.465 ;
        RECT  15.700 3.660 16.115 3.965 ;
        RECT  15.680 0.700 16.070 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.665 3.995 2.030 4.250 ;
        RECT  1.665 3.960 2.010 4.250 ;
        RECT  1.665 3.470 1.895 4.250 ;
        RECT  1.410 3.470 1.895 3.815 ;
        RECT  1.385 3.470 1.895 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.970 2.800 3.655 3.190 ;
        RECT  2.970 2.045 3.200 3.190 ;
        RECT  0.575 2.045 3.200 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.805 2.650 3.190 ;
        RECT  2.310 2.580 2.650 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 1.660 10.105 2.120 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.310 2.045 14.040 2.580 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.460 1.930 15.090 2.580 ;
        END
    END SN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.005 ;
        RECT  14.385 -0.400 14.725 1.025 ;
        RECT  9.450 -0.400 9.755 0.970 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.390 3.330 16.730 5.280 ;
        RECT  15.085 4.170 15.425 5.280 ;
        RECT  13.295 3.665 13.635 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.855 3.845 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.720 1.815 ;
        RECT  3.380 1.555 3.720 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.310 1.630 ;
        RECT  4.140 1.550 4.480 2.090 ;
        RECT  3.950 1.860 6.710 2.090 ;
        RECT  6.370 1.860 6.710 2.460 ;
        RECT  3.950 1.860 4.180 3.135 ;
        RECT  3.930 2.795 4.270 3.135 ;
        RECT  6.955 1.200 7.540 1.540 ;
        RECT  4.420 2.320 5.535 2.605 ;
        RECT  5.305 2.320 5.535 3.155 ;
        RECT  6.955 1.200 7.185 3.385 ;
        RECT  5.305 2.870 7.185 3.155 ;
        RECT  6.955 3.045 7.510 3.385 ;
        RECT  4.380 3.385 6.725 3.615 ;
        RECT  2.125 3.420 4.505 3.650 ;
        RECT  2.125 3.420 2.410 3.760 ;
        RECT  7.930 3.535 8.270 3.845 ;
        RECT  6.495 3.615 8.270 3.845 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.740 8.230 0.970 ;
        RECT  1.255 1.585 2.30 1.815 ;
        RECT  2.825 1.090 3.40 1.320 ;
        RECT  3.950 1.860 5.60 2.090 ;
        RECT  4.380 3.385 5.50 3.615 ;
        RECT  2.125 3.420 3.20 3.650 ;
        RECT  2.255 0.630 4.60 0.860 ;
        RECT  6.145 0.740 7.40 0.970 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  8.000 0.740 8.230 1.600 ;
        RECT  8.000 1.260 8.340 1.600 ;
        RECT  7.415 1.795 7.700 2.700 ;
        RECT  10.445 1.240 10.675 3.120 ;
        RECT  7.415 2.470 7.970 2.700 ;
        RECT  9.115 2.625 10.675 2.965 ;
        RECT  7.740 2.470 7.970 3.305 ;
        RECT  10.430 2.890 11.785 3.120 ;
        RECT  11.445 2.890 11.785 3.230 ;
        RECT  9.115 2.020 9.345 3.305 ;
        RECT  7.740 3.075 9.345 3.305 ;
        RECT  9.985 0.780 11.135 1.010 ;
        RECT  8.650 0.630 8.990 1.430 ;
        RECT  9.985 0.780 10.215 1.430 ;
        RECT  8.650 1.200 10.215 1.430 ;
        RECT  10.905 0.780 11.135 2.450 ;
        RECT  8.650 0.630 8.885 2.235 ;
        RECT  8.150 1.950 8.770 2.290 ;
        RECT  10.905 2.220 11.655 2.450 ;
        RECT  11.315 2.330 12.420 2.560 ;
        RECT  8.430 1.950 8.770 2.845 ;
        RECT  12.135 2.330 12.420 3.450 ;
        RECT  11.365 0.630 13.960 0.860 ;
        RECT  11.365 0.630 11.650 1.005 ;
        RECT  13.620 0.630 13.960 1.200 ;
        RECT  12.320 1.090 12.880 1.400 ;
        RECT  12.650 2.810 15.145 3.040 ;
        RECT  12.650 2.810 14.170 3.070 ;
        RECT  12.650 1.090 12.880 3.970 ;
        RECT  11.725 3.680 12.880 3.970 ;
        RECT  13.270 1.425 13.570 1.740 ;
        RECT  13.270 1.435 15.605 1.665 ;
        RECT  13.270 1.435 13.610 1.740 ;
        RECT  15.375 1.695 15.920 1.980 ;
        RECT  15.375 2.300 16.170 2.640 ;
        RECT  15.375 1.435 15.605 3.450 ;
        RECT  14.285 3.270 15.525 3.500 ;
        RECT  14.285 3.270 14.625 4.005 ;
    END
END SDFRRSX1

MACRO SDFRRSX0
    CLASS CORE ;
    FOREIGN SDFRRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.305 3.810 16.885 4.165 ;
        RECT  16.485 2.860 16.885 4.165 ;
        RECT  16.485 1.170 16.715 4.165 ;
        RECT  16.265 1.170 16.715 1.500 ;
        RECT  16.255 1.170 16.715 1.455 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.455  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.395 2.550 16.070 2.780 ;
        RECT  15.840 1.625 16.070 2.780 ;
        RECT  15.770 0.630 16.000 1.810 ;
        RECT  15.175 0.630 16.000 0.950 ;
        RECT  15.250 2.860 15.625 3.350 ;
        RECT  15.395 2.550 15.625 3.350 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.260 2.415 2.550 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.240 9.665 2.660 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.245 13.350 2.750 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 2.250 14.560 2.680 ;
        END
    END SN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.250 3.810 15.595 5.280 ;
        RECT  12.715 3.910 13.520 5.280 ;
        RECT  9.940 3.630 10.280 5.280 ;
        RECT  8.655 3.940 8.995 5.280 ;
        RECT  4.830 3.865 5.620 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.255 -0.400 16.595 0.710 ;
        RECT  14.145 -0.400 14.485 0.950 ;
        RECT  9.045 -0.400 9.330 1.400 ;
        RECT  4.715 -0.400 5.055 0.710 ;
        RECT  0.180 -0.400 0.520 1.570 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.800 1.320 2.030 ;
        RECT  0.245 1.800 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.500 1.090 3.730 1.630 ;
        RECT  5.565 1.395 5.855 1.630 ;
        RECT  3.500 1.400 5.855 1.630 ;
        RECT  3.505 1.860 5.955 2.120 ;
        RECT  5.670 1.860 5.955 2.205 ;
        RECT  3.505 1.860 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  6.185 1.230 7.085 1.540 ;
        RECT  3.965 2.350 5.275 2.665 ;
        RECT  4.930 2.350 5.275 3.175 ;
        RECT  4.930 2.945 6.415 3.175 ;
        RECT  6.185 1.230 6.415 3.250 ;
        RECT  6.245 3.080 6.825 3.310 ;
        RECT  6.595 3.080 6.825 3.790 ;
        RECT  6.595 3.450 6.935 3.790 ;
        RECT  4.370 3.450 6.040 3.635 ;
        RECT  4.370 3.405 6.010 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.850 3.475 6.080 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.355 3.940 7.695 4.250 ;
        RECT  5.850 4.020 7.695 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  3.960 0.630 4.190 1.170 ;
        RECT  5.285 0.770 7.885 1.000 ;
        RECT  3.960 0.940 5.515 1.170 ;
        RECT  7.545 0.770 7.885 1.570 ;
        RECT  8.305 2.395 8.655 2.735 ;
        RECT  6.645 2.510 7.395 2.850 ;
        RECT  10.020 1.230 10.250 3.360 ;
        RECT  10.020 3.020 11.230 3.360 ;
        RECT  8.425 3.110 11.230 3.360 ;
        RECT  8.425 3.110 9.595 3.450 ;
        RECT  7.165 2.510 7.395 3.710 ;
        RECT  8.425 2.395 8.655 3.710 ;
        RECT  7.165 3.480 8.655 3.710 ;
        RECT  9.560 0.770 10.710 1.000 ;
        RECT  8.245 1.230 8.585 1.870 ;
        RECT  8.245 1.640 9.790 1.870 ;
        RECT  9.560 0.770 9.790 1.870 ;
        RECT  10.480 0.770 10.710 2.290 ;
        RECT  6.645 1.840 8.475 2.110 ;
        RECT  6.645 1.840 8.075 2.180 ;
        RECT  10.480 2.060 11.245 2.290 ;
        RECT  10.905 2.170 11.915 2.400 ;
        RECT  7.845 1.840 8.075 3.250 ;
        RECT  11.685 2.170 11.915 3.440 ;
        RECT  7.845 2.965 8.195 3.250 ;
        RECT  11.685 3.100 12.025 3.440 ;
        RECT  10.940 0.630 13.685 0.860 ;
        RECT  13.345 0.630 13.685 1.200 ;
        RECT  10.940 0.630 11.225 1.400 ;
        RECT  12.115 1.090 12.485 1.400 ;
        RECT  12.255 3.125 14.525 3.465 ;
        RECT  12.255 1.090 12.485 3.970 ;
        RECT  11.235 3.670 12.485 3.970 ;
        RECT  13.075 1.430 15.515 1.775 ;
        RECT  15.175 1.350 15.515 2.320 ;
        RECT  14.790 1.430 15.515 2.320 ;
        RECT  14.790 1.980 15.610 2.320 ;
        RECT  14.790 1.430 15.020 4.175 ;
        RECT  14.205 3.835 15.020 4.175 ;
        RECT  0.980 1.585 2.80 1.960 ;
        RECT  1.445 1.125 2.80 1.355 ;
        RECT  3.500 1.400 4.70 1.630 ;
        RECT  3.505 1.860 4.00 2.120 ;
        RECT  1.995 3.710 3.60 3.940 ;
        RECT  1.980 0.630 3.50 0.860 ;
        RECT  5.285 0.770 6.60 1.000 ;
        RECT  8.425 3.110 10.60 3.360 ;
        RECT  10.940 0.630 12.30 0.860 ;
        RECT  12.255 3.125 13.20 3.465 ;
        RECT  13.075 1.430 14.40 1.775 ;
    END
END SDFRRSX0

MACRO SDFRRSQX4
    CLASS CORE ;
    FOREIGN SDFRRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 1.130 19.980 4.030 ;
        RECT  18.200 2.250 19.980 2.630 ;
        RECT  18.200 1.130 18.540 4.030 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.875 1.640 16.365 2.150 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.175 2.180 15.645 2.700 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 1.660 11.015 2.100 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.470 ;
        RECT  17.440 -0.400 17.780 0.800 ;
        RECT  15.875 -0.400 16.215 0.760 ;
        RECT  10.350 -0.400 10.635 0.970 ;
        RECT  4.775 -0.400 6.345 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  18.920 2.860 19.260 5.280 ;
        RECT  17.440 4.070 17.780 5.280 ;
        RECT  14.955 3.910 16.415 5.280 ;
        RECT  12.655 3.965 12.995 5.280 ;
        RECT  10.235 2.910 10.535 5.280 ;
        RECT  4.830 3.965 6.300 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 6.485 2.095 ;
        RECT  6.255 1.860 6.485 2.800 ;
        RECT  6.255 2.460 6.595 2.800 ;
        RECT  3.895 1.815 4.125 3.370 ;
        RECT  3.895 3.085 4.260 3.370 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 7.055 1.585 ;
        RECT  5.445 1.355 7.055 1.630 ;
        RECT  6.765 1.355 7.055 1.695 ;
        RECT  7.285 1.160 8.330 1.500 ;
        RECT  4.355 2.325 4.640 2.665 ;
        RECT  4.355 2.435 5.490 2.665 ;
        RECT  5.260 2.435 5.490 3.275 ;
        RECT  5.260 2.935 5.600 3.275 ;
        RECT  7.285 1.160 7.515 3.540 ;
        RECT  5.260 3.045 7.515 3.275 ;
        RECT  7.200 3.200 7.545 3.540 ;
        RECT  4.450 3.505 6.820 3.735 ;
        RECT  6.590 3.505 6.820 4.000 ;
        RECT  2.020 3.600 4.640 3.830 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  8.010 2.980 8.350 4.000 ;
        RECT  6.590 3.770 8.350 4.000 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.640 0.700 8.790 0.930 ;
        RECT  4.315 0.895 6.870 1.125 ;
        RECT  8.560 0.700 8.790 1.660 ;
        RECT  8.560 1.320 9.145 1.660 ;
        RECT  10.865 0.775 12.015 1.005 ;
        RECT  9.020 0.735 9.890 1.090 ;
        RECT  10.865 0.775 11.095 1.430 ;
        RECT  9.660 1.200 11.095 1.430 ;
        RECT  11.785 0.775 12.015 2.090 ;
        RECT  11.785 1.860 13.450 2.090 ;
        RECT  9.660 0.735 9.890 2.150 ;
        RECT  9.260 1.920 9.890 2.150 ;
        RECT  13.110 1.860 13.450 2.200 ;
        RECT  9.260 1.920 9.545 3.195 ;
        RECT  7.745 1.890 9.030 2.120 ;
        RECT  7.745 1.810 8.055 2.175 ;
        RECT  11.325 1.240 11.555 2.680 ;
        RECT  11.325 2.340 12.025 2.680 ;
        RECT  13.780 1.670 14.065 2.680 ;
        RECT  9.775 2.450 14.065 2.680 ;
        RECT  10.915 2.450 11.255 2.860 ;
        RECT  8.690 1.890 9.030 3.655 ;
        RECT  10.915 2.450 11.145 3.855 ;
        RECT  9.775 2.450 10.005 3.655 ;
        RECT  8.690 3.425 10.005 3.655 ;
        RECT  12.125 3.505 13.635 3.735 ;
        RECT  13.405 3.505 13.635 4.100 ;
        RECT  10.915 3.625 12.355 3.855 ;
        RECT  13.405 3.760 13.745 4.100 ;
        RECT  12.245 0.630 15.210 0.860 ;
        RECT  14.870 0.630 15.210 0.950 ;
        RECT  12.245 0.630 12.540 1.500 ;
        RECT  13.350 1.100 13.690 1.440 ;
        RECT  13.350 1.210 14.525 1.440 ;
        RECT  17.025 2.270 17.365 2.610 ;
        RECT  16.375 2.380 17.365 2.610 ;
        RECT  14.295 1.210 14.525 3.275 ;
        RECT  16.375 2.380 16.605 3.275 ;
        RECT  11.465 3.045 16.605 3.275 ;
        RECT  15.515 3.045 15.855 3.385 ;
        RECT  11.465 3.045 11.805 3.395 ;
        RECT  13.975 3.045 14.265 3.780 ;
        RECT  14.755 1.180 17.280 1.410 ;
        RECT  16.940 1.350 17.825 1.580 ;
        RECT  14.755 1.180 15.095 1.675 ;
        RECT  17.595 1.350 17.825 3.070 ;
        RECT  16.835 2.840 17.825 3.070 ;
        RECT  16.835 2.840 17.175 3.660 ;
        RECT  1.145 1.585 2.80 1.815 ;
        RECT  3.895 1.860 5.40 2.095 ;
        RECT  1.605 1.125 3.90 1.355 ;
        RECT  3.855 1.355 6.50 1.585 ;
        RECT  5.260 3.045 6.60 3.275 ;
        RECT  4.450 3.505 5.80 3.735 ;
        RECT  2.020 3.600 3.50 3.830 ;
        RECT  2.255 0.630 3.70 0.895 ;
        RECT  6.640 0.700 7.70 0.930 ;
        RECT  4.315 0.895 5.30 1.125 ;
        RECT  9.775 2.450 13.20 2.680 ;
        RECT  12.245 0.630 14.60 0.860 ;
        RECT  11.465 3.045 15.80 3.275 ;
        RECT  14.755 1.180 16.90 1.410 ;
    END
END SDFRRSQX4

MACRO SDFRRSQX2
    CLASS CORE ;
    FOREIGN SDFRRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.560 1.240 16.900 2.630 ;
        RECT  16.340 2.250 16.735 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.020 10.040 2.630 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 2.035 14.125 2.375 ;
        RECT  13.355 2.035 13.735 2.630 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.050 14.995 2.630 ;
        RECT  14.475 2.050 14.995 2.395 ;
        END
    END SN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  17.120 -0.400 17.460 0.720 ;
        RECT  16.000 -0.400 16.340 0.720 ;
        RECT  14.395 -0.400 14.735 0.970 ;
        RECT  9.385 -0.400 9.670 1.330 ;
        RECT  5.630 -0.400 5.920 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  17.060 3.270 17.400 5.280 ;
        RECT  15.580 4.170 15.920 5.280 ;
        RECT  14.260 3.910 14.600 5.280 ;
        RECT  13.120 3.825 13.460 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.965 3.900 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.265 1.630 ;
        RECT  4.135 1.550 4.475 2.090 ;
        RECT  3.895 1.860 6.545 2.090 ;
        RECT  6.205 1.860 6.545 2.375 ;
        RECT  3.895 1.860 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.850 1.190 7.495 1.530 ;
        RECT  4.355 2.320 5.645 2.635 ;
        RECT  6.850 1.190 7.080 3.210 ;
        RECT  5.305 2.320 5.645 3.210 ;
        RECT  6.850 2.870 7.510 3.210 ;
        RECT  5.305 2.980 7.510 3.210 ;
        RECT  4.505 3.440 6.705 3.670 ;
        RECT  2.120 3.500 4.735 3.730 ;
        RECT  7.930 3.535 8.270 3.845 ;
        RECT  6.475 3.615 8.270 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.150 0.730 8.295 0.960 ;
        RECT  5.170 0.940 6.380 1.170 ;
        RECT  7.955 0.730 8.295 1.600 ;
        RECT  9.900 0.800 11.050 1.030 ;
        RECT  8.570 0.630 8.950 1.790 ;
        RECT  10.820 0.800 11.050 1.790 ;
        RECT  9.900 0.800 10.130 1.790 ;
        RECT  8.570 1.560 10.130 1.790 ;
        RECT  10.820 1.560 12.475 1.790 ;
        RECT  12.135 1.560 12.475 1.895 ;
        RECT  8.240 2.020 8.800 2.360 ;
        RECT  8.570 0.630 8.800 2.845 ;
        RECT  8.460 2.020 8.800 2.845 ;
        RECT  7.310 1.795 7.650 2.115 ;
        RECT  7.310 1.885 7.970 2.115 ;
        RECT  11.245 2.120 11.585 2.460 ;
        RECT  11.245 2.225 12.630 2.460 ;
        RECT  10.360 2.230 12.630 2.460 ;
        RECT  12.345 2.225 12.630 2.565 ;
        RECT  9.030 2.020 9.345 3.145 ;
        RECT  7.740 1.885 7.970 3.305 ;
        RECT  9.030 2.860 10.590 3.145 ;
        RECT  10.360 1.260 10.590 3.145 ;
        RECT  7.740 3.075 9.260 3.305 ;
        RECT  11.280 0.630 13.975 0.860 ;
        RECT  13.635 0.630 13.975 1.105 ;
        RECT  11.280 0.630 11.565 1.330 ;
        RECT  12.405 1.090 13.090 1.330 ;
        RECT  12.860 1.090 13.090 3.090 ;
        RECT  13.965 2.605 14.305 3.090 ;
        RECT  15.225 2.750 15.565 3.090 ;
        RECT  11.725 2.860 15.565 3.090 ;
        RECT  11.725 2.860 12.065 3.615 ;
        RECT  15.225 0.630 15.565 1.610 ;
        RECT  13.355 1.380 16.025 1.610 ;
        RECT  13.355 1.380 13.700 1.720 ;
        RECT  15.795 1.380 16.025 3.610 ;
        RECT  15.020 3.380 16.025 3.610 ;
        RECT  15.020 3.380 15.360 3.720 ;
        RECT  1.255 1.585 2.50 1.815 ;
        RECT  2.825 1.090 3.60 1.320 ;
        RECT  1.715 1.125 2.70 1.355 ;
        RECT  3.895 1.860 5.60 2.090 ;
        RECT  5.305 2.980 6.90 3.210 ;
        RECT  4.505 3.440 5.70 3.670 ;
        RECT  2.120 3.500 3.60 3.730 ;
        RECT  2.255 0.630 4.70 0.860 ;
        RECT  6.150 0.730 7.60 0.960 ;
        RECT  10.360 2.230 11.80 2.460 ;
        RECT  11.280 0.630 12.30 0.860 ;
        RECT  11.725 2.860 14.40 3.090 ;
        RECT  13.355 1.380 15.60 1.610 ;
    END
END SDFRRSQX2

MACRO SDFRRSQX1
    CLASS CORE ;
    FOREIGN SDFRRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.875 2.250 16.380 2.635 ;
        RECT  16.150 1.235 16.380 2.635 ;
        RECT  15.840 1.235 16.380 1.465 ;
        RECT  15.670 3.680 16.115 3.965 ;
        RECT  15.875 2.250 16.115 3.965 ;
        RECT  15.840 0.700 16.070 1.465 ;
        RECT  15.700 3.660 16.115 3.965 ;
        RECT  15.680 0.700 16.070 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.665 3.995 2.030 4.250 ;
        RECT  1.665 3.960 2.010 4.250 ;
        RECT  1.665 3.470 1.895 4.250 ;
        RECT  1.410 3.470 1.895 3.815 ;
        RECT  1.385 3.470 1.895 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.970 2.800 3.655 3.190 ;
        RECT  2.970 2.045 3.200 3.190 ;
        RECT  0.575 2.045 3.200 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 1.660 10.105 2.120 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.310 2.045 14.040 2.580 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.460 1.930 15.090 2.580 ;
        END
    END SN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.400 -0.400 16.740 1.005 ;
        RECT  14.385 -0.400 14.725 1.025 ;
        RECT  9.450 -0.400 9.755 0.970 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.390 3.330 16.730 5.280 ;
        RECT  15.085 4.170 15.425 5.280 ;
        RECT  13.295 3.665 13.635 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.855 3.845 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.720 1.815 ;
        RECT  3.380 1.555 3.720 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.310 1.630 ;
        RECT  4.140 1.550 4.480 2.090 ;
        RECT  3.950 1.860 6.710 2.090 ;
        RECT  6.370 1.860 6.710 2.460 ;
        RECT  3.950 1.860 4.180 3.135 ;
        RECT  3.930 2.795 4.270 3.135 ;
        RECT  6.955 1.200 7.540 1.540 ;
        RECT  4.420 2.320 5.535 2.605 ;
        RECT  5.305 2.320 5.535 3.155 ;
        RECT  6.955 1.200 7.185 3.385 ;
        RECT  5.305 2.870 7.185 3.155 ;
        RECT  6.955 3.045 7.510 3.385 ;
        RECT  4.380 3.385 6.725 3.615 ;
        RECT  2.125 3.420 4.505 3.650 ;
        RECT  2.125 3.420 2.410 3.760 ;
        RECT  7.930 3.535 8.270 3.845 ;
        RECT  6.495 3.615 8.270 3.845 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.740 8.230 0.970 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  8.000 0.740 8.230 1.600 ;
        RECT  8.000 1.260 8.340 1.600 ;
        RECT  7.415 1.800 7.700 2.700 ;
        RECT  10.445 1.240 10.675 3.120 ;
        RECT  7.415 2.470 7.970 2.700 ;
        RECT  9.115 2.625 10.675 2.965 ;
        RECT  7.740 2.470 7.970 3.305 ;
        RECT  10.430 2.890 11.785 3.120 ;
        RECT  11.445 2.890 11.785 3.230 ;
        RECT  9.115 2.020 9.345 3.305 ;
        RECT  7.740 3.075 9.345 3.305 ;
        RECT  9.985 0.780 11.135 1.010 ;
        RECT  8.650 0.630 8.990 1.430 ;
        RECT  9.985 0.780 10.215 1.430 ;
        RECT  8.650 1.200 10.215 1.430 ;
        RECT  10.905 0.780 11.135 2.450 ;
        RECT  8.650 0.630 8.885 2.235 ;
        RECT  8.150 1.950 8.770 2.290 ;
        RECT  10.905 2.220 11.655 2.450 ;
        RECT  11.315 2.330 12.420 2.560 ;
        RECT  8.430 1.950 8.770 2.845 ;
        RECT  12.135 2.330 12.420 3.450 ;
        RECT  11.365 0.630 13.960 0.860 ;
        RECT  11.365 0.630 11.650 1.005 ;
        RECT  13.620 0.630 13.960 1.200 ;
        RECT  12.320 1.090 12.880 1.400 ;
        RECT  12.650 2.810 15.145 3.040 ;
        RECT  12.650 2.810 14.170 3.070 ;
        RECT  12.650 1.090 12.880 3.970 ;
        RECT  11.725 3.680 12.880 3.970 ;
        RECT  13.270 1.425 13.570 1.740 ;
        RECT  13.270 1.435 15.605 1.665 ;
        RECT  13.270 1.435 13.610 1.740 ;
        RECT  15.375 1.695 15.920 1.980 ;
        RECT  15.375 1.435 15.605 3.450 ;
        RECT  14.285 3.270 15.525 3.500 ;
        RECT  14.285 3.270 14.625 4.005 ;
        RECT  1.255 1.585 2.70 1.815 ;
        RECT  2.825 1.090 3.60 1.320 ;
        RECT  3.950 1.860 5.60 2.090 ;
        RECT  4.380 3.385 5.90 3.615 ;
        RECT  2.125 3.420 3.70 3.650 ;
        RECT  2.255 0.630 4.00 0.860 ;
        RECT  6.145 0.740 7.30 0.970 ;
        RECT  11.365 0.630 12.20 0.860 ;
        RECT  12.650 2.810 14.70 3.040 ;
        RECT  13.270 1.435 14.70 1.665 ;
    END
END SDFRRSQX1

MACRO SDFRRSQX0
    CLASS CORE ;
    FOREIGN SDFRRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.512  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.220 2.860 15.635 3.350 ;
        RECT  15.405 0.635 15.635 3.350 ;
        RECT  14.855 0.635 15.635 0.975 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.260 2.415 2.550 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.240 9.665 2.660 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.250 13.380 2.895 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 2.285 14.485 2.795 ;
        END
    END SN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.220 3.810 15.560 5.280 ;
        RECT  12.715 3.910 13.520 5.280 ;
        RECT  9.940 3.630 10.280 5.280 ;
        RECT  8.655 3.940 8.995 5.280 ;
        RECT  4.830 3.865 5.620 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  13.825 -0.400 14.165 0.975 ;
        RECT  9.045 -0.400 9.330 1.400 ;
        RECT  4.715 -0.400 5.055 0.710 ;
        RECT  0.180 -0.400 0.520 1.570 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.800 1.320 2.030 ;
        RECT  0.245 1.800 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.500 1.090 3.730 1.630 ;
        RECT  5.565 1.395 5.855 1.630 ;
        RECT  3.500 1.400 5.855 1.630 ;
        RECT  3.505 1.860 5.950 2.120 ;
        RECT  5.665 1.860 5.950 2.205 ;
        RECT  3.505 1.860 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  6.180 1.230 7.085 1.540 ;
        RECT  3.965 2.350 5.275 2.665 ;
        RECT  4.930 2.350 5.275 3.175 ;
        RECT  4.930 2.945 6.410 3.175 ;
        RECT  6.180 1.230 6.410 3.175 ;
        RECT  6.235 3.025 6.825 3.255 ;
        RECT  6.595 3.025 6.825 3.790 ;
        RECT  6.595 3.450 6.935 3.790 ;
        RECT  4.370 3.405 6.055 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.850 3.435 6.080 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.355 3.940 7.695 4.250 ;
        RECT  5.850 4.020 7.695 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  3.960 0.630 4.190 1.170 ;
        RECT  5.285 0.770 7.885 1.000 ;
        RECT  3.960 0.940 5.515 1.170 ;
        RECT  7.545 0.770 7.885 1.570 ;
        RECT  6.640 2.510 6.975 2.795 ;
        RECT  8.305 2.395 8.655 2.735 ;
        RECT  6.640 2.530 7.395 2.795 ;
        RECT  10.020 1.230 10.250 3.395 ;
        RECT  10.020 3.055 11.230 3.395 ;
        RECT  8.425 3.110 11.230 3.395 ;
        RECT  8.425 3.110 9.595 3.450 ;
        RECT  7.165 2.530 7.395 3.710 ;
        RECT  8.425 2.395 8.655 3.710 ;
        RECT  7.165 3.480 8.655 3.710 ;
        RECT  9.560 0.770 10.710 1.000 ;
        RECT  8.245 1.230 8.585 1.870 ;
        RECT  8.245 1.640 9.790 1.870 ;
        RECT  9.560 0.770 9.790 1.870 ;
        RECT  6.640 1.840 8.475 2.110 ;
        RECT  6.640 1.840 8.075 2.180 ;
        RECT  10.480 0.770 10.710 2.480 ;
        RECT  10.480 2.235 12.025 2.480 ;
        RECT  7.845 1.840 8.075 3.250 ;
        RECT  7.845 2.965 8.195 3.250 ;
        RECT  11.685 2.235 12.025 3.440 ;
        RECT  10.940 0.635 13.280 0.865 ;
        RECT  10.940 0.635 11.225 0.975 ;
        RECT  12.940 0.635 13.280 0.975 ;
        RECT  11.915 1.175 12.485 1.515 ;
        RECT  13.235 3.125 14.525 3.465 ;
        RECT  12.255 3.235 14.525 3.465 ;
        RECT  12.255 1.175 12.485 3.970 ;
        RECT  11.235 3.670 12.485 3.970 ;
        RECT  14.760 1.350 15.175 1.690 ;
        RECT  12.875 1.735 14.990 2.020 ;
        RECT  14.760 1.350 14.990 4.175 ;
        RECT  14.160 3.835 14.990 4.175 ;
        RECT  0.980 1.585 2.60 1.960 ;
        RECT  1.445 1.125 2.50 1.355 ;
        RECT  3.500 1.400 4.80 1.630 ;
        RECT  3.505 1.860 4.20 2.120 ;
        RECT  1.995 3.710 3.30 3.940 ;
        RECT  1.980 0.630 3.20 0.860 ;
        RECT  5.285 0.770 6.50 1.000 ;
        RECT  8.425 3.110 10.10 3.395 ;
        RECT  10.940 0.635 12.40 0.865 ;
        RECT  12.255 3.235 13.80 3.465 ;
        RECT  12.875 1.735 13.40 2.020 ;
    END
END SDFRRSQX0

MACRO SDFRRQX4
    CLASS CORE ;
    FOREIGN SDFRRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.010 1.130 19.350 4.010 ;
        RECT  17.570 2.250 19.350 2.630 ;
        RECT  17.570 1.130 17.910 4.010 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.020 1.640 15.625 2.100 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.660 10.630 2.135 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.290 -0.400 18.630 1.470 ;
        RECT  16.810 -0.400 17.150 0.725 ;
        RECT  15.500 -0.400 15.840 0.950 ;
        RECT  9.920 -0.400 10.205 0.970 ;
        RECT  4.775 -0.400 5.915 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.290 2.860 18.630 5.280 ;
        RECT  16.850 2.770 17.190 5.280 ;
        RECT  14.155 3.760 15.615 5.280 ;
        RECT  12.095 3.980 12.435 5.280 ;
        RECT  9.540 2.950 9.825 5.280 ;
        RECT  4.660 4.115 5.700 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 5.885 2.095 ;
        RECT  5.655 1.860 5.885 2.800 ;
        RECT  5.655 2.460 5.995 2.800 ;
        RECT  3.895 1.815 4.125 3.425 ;
        RECT  3.895 3.085 4.260 3.425 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 6.625 1.585 ;
        RECT  5.015 1.355 6.625 1.630 ;
        RECT  6.335 1.355 6.625 1.695 ;
        RECT  2.020 3.655 6.390 3.885 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  6.160 3.850 7.710 4.080 ;
        RECT  7.370 3.850 7.710 4.190 ;
        RECT  6.855 1.160 7.900 1.500 ;
        RECT  4.355 2.325 4.640 2.665 ;
        RECT  4.355 2.435 4.890 2.665 ;
        RECT  4.660 2.435 4.890 3.425 ;
        RECT  4.660 3.085 5.000 3.425 ;
        RECT  4.660 3.195 7.085 3.425 ;
        RECT  6.855 1.160 7.085 3.540 ;
        RECT  6.745 3.195 7.085 3.540 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.210 0.700 8.360 0.930 ;
        RECT  4.315 0.895 6.440 1.125 ;
        RECT  8.130 0.700 8.360 1.660 ;
        RECT  8.130 1.320 8.715 1.660 ;
        RECT  10.435 0.775 11.585 1.005 ;
        RECT  8.590 0.735 9.460 1.090 ;
        RECT  10.435 0.775 10.665 1.430 ;
        RECT  9.230 1.200 10.665 1.430 ;
        RECT  11.355 0.775 11.585 2.090 ;
        RECT  11.355 1.860 13.020 2.090 ;
        RECT  9.230 0.735 9.460 2.150 ;
        RECT  8.620 1.920 9.460 2.150 ;
        RECT  12.680 1.860 13.020 2.200 ;
        RECT  8.620 1.920 8.850 3.580 ;
        RECT  8.510 3.235 8.850 3.580 ;
        RECT  13.350 1.670 13.690 2.010 ;
        RECT  7.315 1.805 7.625 2.175 ;
        RECT  10.895 1.240 11.125 2.680 ;
        RECT  10.895 2.340 11.485 2.680 ;
        RECT  13.350 1.670 13.580 2.680 ;
        RECT  9.080 2.450 13.580 2.680 ;
        RECT  7.395 1.805 7.625 3.095 ;
        RECT  7.395 2.865 8.280 3.095 ;
        RECT  7.940 2.865 8.280 3.205 ;
        RECT  10.205 2.450 10.545 3.915 ;
        RECT  11.565 3.520 12.895 3.750 ;
        RECT  8.050 2.865 8.280 4.040 ;
        RECT  12.665 3.520 12.895 4.200 ;
        RECT  10.205 3.685 11.795 3.915 ;
        RECT  9.080 2.450 9.310 4.040 ;
        RECT  8.050 3.810 9.310 4.040 ;
        RECT  12.665 3.860 13.185 4.200 ;
        RECT  11.815 0.630 15.040 0.860 ;
        RECT  14.230 0.630 15.040 0.950 ;
        RECT  11.815 0.630 12.110 1.500 ;
        RECT  12.920 1.090 13.260 1.440 ;
        RECT  12.920 1.210 14.150 1.440 ;
        RECT  15.800 2.250 16.140 2.590 ;
        RECT  13.920 2.360 16.140 2.590 ;
        RECT  14.715 2.360 15.055 3.150 ;
        RECT  13.920 1.210 14.150 3.215 ;
        RECT  10.905 2.985 14.150 3.215 ;
        RECT  10.905 2.985 11.245 3.455 ;
        RECT  13.125 2.985 13.465 3.630 ;
        RECT  14.380 1.180 16.600 1.410 ;
        RECT  16.260 1.080 16.600 1.420 ;
        RECT  14.380 1.180 14.720 1.675 ;
        RECT  16.370 1.080 16.600 3.640 ;
        RECT  16.130 2.820 16.600 3.640 ;
        RECT  1.145 1.585 2.40 1.815 ;
        RECT  1.605 1.125 3.30 1.355 ;
        RECT  3.855 1.355 5.20 1.585 ;
        RECT  2.020 3.655 5.50 3.885 ;
        RECT  4.660 3.195 6.00 3.425 ;
        RECT  2.255 0.630 3.40 0.895 ;
        RECT  6.210 0.700 7.80 0.930 ;
        RECT  4.315 0.895 5.40 1.125 ;
        RECT  9.080 2.450 12.90 2.680 ;
        RECT  11.815 0.630 14.40 0.860 ;
        RECT  13.920 2.360 15.90 2.590 ;
        RECT  10.905 2.985 13.30 3.215 ;
        RECT  14.380 1.180 15.20 1.410 ;
    END
END SDFRRQX4

MACRO SDFRRQX2
    CLASS CORE ;
    FOREIGN SDFRRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.020 0.820 16.255 3.240 ;
        RECT  15.770 2.860 16.110 3.830 ;
        RECT  15.770 0.820 16.255 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.250 9.700 2.630 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.200 2.110 13.735 2.675 ;
        END
    END RN
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 1.160 ;
        RECT  15.050 -0.400 15.390 1.160 ;
        RECT  14.005 -0.400 14.345 1.220 ;
        RECT  9.035 -0.400 9.320 1.330 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.490 2.920 16.830 5.280 ;
        RECT  15.010 3.775 15.350 5.280 ;
        RECT  12.745 3.365 13.085 5.280 ;
        RECT  9.895 3.525 10.235 5.280 ;
        RECT  8.595 3.810 8.935 5.280 ;
        RECT  4.655 3.960 5.645 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.685 ;
        RECT  4.710 1.400 5.915 1.685 ;
        RECT  4.135 1.550 4.475 2.180 ;
        RECT  3.895 1.950 6.165 2.180 ;
        RECT  5.825 1.950 6.165 2.375 ;
        RECT  3.895 1.950 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.805 1.260 7.145 1.600 ;
        RECT  6.495 1.370 7.145 1.600 ;
        RECT  4.415 2.410 5.045 2.750 ;
        RECT  4.705 2.410 5.045 3.270 ;
        RECT  6.495 1.370 6.725 3.270 ;
        RECT  4.705 3.040 6.875 3.270 ;
        RECT  6.535 3.040 6.875 3.625 ;
        RECT  2.120 3.500 6.305 3.730 ;
        RECT  6.075 3.500 6.305 4.125 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  7.295 3.810 7.635 4.125 ;
        RECT  6.075 3.895 7.635 4.125 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.800 7.945 1.030 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  7.605 0.800 7.945 1.600 ;
        RECT  9.550 0.800 10.700 1.030 ;
        RECT  8.260 0.630 8.600 1.790 ;
        RECT  10.470 0.800 10.700 1.790 ;
        RECT  9.550 0.800 9.780 1.790 ;
        RECT  8.260 1.560 9.780 1.790 ;
        RECT  10.470 1.560 12.125 1.790 ;
        RECT  11.785 1.560 12.125 1.895 ;
        RECT  8.260 0.630 8.490 2.060 ;
        RECT  7.755 1.830 8.490 2.060 ;
        RECT  7.755 1.830 8.165 2.240 ;
        RECT  7.825 1.830 8.165 3.120 ;
        RECT  6.955 1.900 7.335 2.215 ;
        RECT  10.810 2.225 12.320 2.565 ;
        RECT  10.010 2.230 12.320 2.565 ;
        RECT  8.425 2.305 8.715 3.165 ;
        RECT  10.010 1.260 10.240 3.165 ;
        RECT  8.425 2.860 10.240 3.165 ;
        RECT  7.105 1.900 7.335 3.580 ;
        RECT  8.425 2.305 8.670 3.580 ;
        RECT  7.105 3.350 8.670 3.580 ;
        RECT  10.930 0.630 13.625 0.860 ;
        RECT  13.285 0.630 13.625 1.105 ;
        RECT  10.930 0.630 11.215 1.330 ;
        RECT  12.055 1.090 12.780 1.330 ;
        RECT  13.965 2.400 14.935 2.740 ;
        RECT  12.550 1.090 12.780 3.135 ;
        RECT  13.965 2.400 14.195 3.135 ;
        RECT  11.300 2.905 14.195 3.135 ;
        RECT  11.300 2.905 11.640 3.690 ;
        RECT  13.465 2.905 13.805 4.175 ;
        RECT  13.010 1.380 13.355 1.720 ;
        RECT  13.010 1.490 15.145 1.720 ;
        RECT  14.805 1.490 15.145 1.980 ;
        RECT  14.805 1.750 15.395 1.980 ;
        RECT  15.165 1.750 15.395 3.200 ;
        RECT  14.450 2.970 15.395 3.200 ;
        RECT  14.450 2.970 14.790 3.310 ;
        RECT  1.255 1.585 2.80 1.815 ;
        RECT  2.825 1.090 3.60 1.320 ;
        RECT  1.715 1.125 2.30 1.355 ;
        RECT  3.895 1.950 5.20 2.180 ;
        RECT  4.705 3.040 5.50 3.270 ;
        RECT  2.120 3.500 5.00 3.730 ;
        RECT  2.255 0.630 4.40 0.860 ;
        RECT  10.010 2.230 11.60 2.565 ;
        RECT  10.930 0.630 12.50 0.860 ;
        RECT  11.300 2.905 13.10 3.135 ;
        RECT  13.010 1.490 14.40 1.720 ;
    END
END SDFRRQX2

MACRO SDFRRQX1
    CLASS CORE ;
    FOREIGN SDFRRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.735 2.250 15.635 2.630 ;
        RECT  14.735 2.250 14.970 3.100 ;
        RECT  14.420 3.780 14.965 4.065 ;
        RECT  14.735 0.700 14.965 4.065 ;
        RECT  14.505 0.700 14.965 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 3.995 2.030 4.250 ;
        RECT  1.610 3.980 2.000 4.250 ;
        RECT  1.610 3.470 1.840 4.250 ;
        RECT  1.410 3.470 1.840 3.815 ;
        RECT  1.385 3.470 1.840 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.980 2.800 3.655 3.240 ;
        RECT  2.980 2.045 3.210 3.240 ;
        RECT  0.575 2.045 3.210 2.275 ;
        RECT  0.575 1.660 0.860 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.030 1.660 9.480 2.130 ;
        RECT  8.945 1.660 9.480 2.030 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.745 2.170 13.290 2.630 ;
        END
    END RN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.195 3.330 15.535 5.280 ;
        RECT  12.740 3.820 13.085 5.280 ;
        RECT  10.125 3.480 10.465 5.280 ;
        RECT  8.825 3.535 9.165 5.280 ;
        RECT  8.870 3.530 9.165 5.280 ;
        RECT  4.910 3.845 5.870 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.225 -0.400 15.565 1.040 ;
        RECT  13.470 -0.400 13.810 0.950 ;
        RECT  8.820 -0.400 9.105 0.970 ;
        RECT  4.815 -0.400 5.155 0.655 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.130 0.900 1.430 ;
        RECT  0.115 1.185 1.485 1.430 ;
        RECT  1.255 1.185 1.485 1.815 ;
        RECT  1.255 1.585 3.665 1.815 ;
        RECT  3.380 1.555 3.665 1.890 ;
        RECT  3.435 1.555 3.665 1.895 ;
        RECT  0.115 1.130 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.410 4.180 ;
        RECT  0.180 3.270 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.125 1.320 ;
        RECT  3.485 1.090 4.125 1.325 ;
        RECT  3.895 1.090 4.125 1.580 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  3.895 1.345 5.685 1.580 ;
        RECT  5.345 1.345 5.685 1.650 ;
        RECT  3.895 1.810 5.165 2.040 ;
        RECT  4.995 1.880 5.960 2.220 ;
        RECT  3.895 1.810 4.215 3.425 ;
        RECT  6.315 1.230 6.915 1.540 ;
        RECT  4.445 2.325 4.755 3.155 ;
        RECT  6.315 1.230 6.545 3.155 ;
        RECT  4.445 2.870 6.545 3.155 ;
        RECT  4.445 2.925 7.095 3.155 ;
        RECT  6.755 2.925 7.095 3.385 ;
        RECT  2.255 0.630 4.585 0.860 ;
        RECT  4.355 0.630 4.585 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.740 0.770 7.660 1.000 ;
        RECT  4.355 0.885 5.970 1.115 ;
        RECT  7.375 0.770 7.660 1.600 ;
        RECT  2.120 3.420 2.405 3.760 ;
        RECT  4.445 3.385 6.330 3.615 ;
        RECT  2.120 3.530 3.575 3.760 ;
        RECT  7.520 3.535 7.860 3.845 ;
        RECT  6.100 3.615 7.860 3.845 ;
        RECT  4.445 3.385 4.675 3.885 ;
        RECT  3.360 3.655 4.675 3.885 ;
        RECT  8.350 2.020 8.715 2.360 ;
        RECT  8.525 2.225 8.820 2.440 ;
        RECT  6.775 1.790 7.065 2.695 ;
        RECT  9.795 1.240 10.025 3.230 ;
        RECT  6.775 2.465 7.555 2.695 ;
        RECT  8.590 2.625 10.025 2.965 ;
        RECT  7.325 2.465 7.555 3.305 ;
        RECT  9.795 2.890 11.375 3.230 ;
        RECT  8.590 2.225 8.820 3.305 ;
        RECT  7.325 3.075 8.820 3.305 ;
        RECT  9.335 0.780 10.485 1.010 ;
        RECT  8.020 0.630 8.360 1.430 ;
        RECT  9.335 0.780 9.565 1.430 ;
        RECT  7.890 1.200 9.565 1.430 ;
        RECT  7.890 1.200 8.120 2.845 ;
        RECT  7.525 1.830 8.120 2.145 ;
        RECT  10.255 0.780 10.485 2.450 ;
        RECT  10.255 2.220 11.095 2.450 ;
        RECT  10.755 2.330 11.840 2.560 ;
        RECT  7.885 1.830 8.120 2.845 ;
        RECT  7.885 2.590 8.350 2.845 ;
        RECT  7.885 2.605 8.360 2.845 ;
        RECT  11.610 2.330 11.840 3.435 ;
        RECT  11.610 3.110 12.050 3.435 ;
        RECT  10.715 0.630 13.040 0.860 ;
        RECT  10.715 0.630 11.000 1.005 ;
        RECT  12.700 0.630 13.040 1.150 ;
        RECT  11.470 1.090 12.300 1.400 ;
        RECT  12.070 1.090 12.300 2.810 ;
        RECT  12.280 2.580 12.515 3.145 ;
        RECT  13.760 2.730 14.045 3.090 ;
        RECT  12.280 2.860 14.045 3.090 ;
        RECT  12.280 2.860 13.580 3.145 ;
        RECT  12.280 2.580 12.510 3.970 ;
        RECT  11.320 3.665 12.510 3.970 ;
        RECT  12.530 1.380 12.815 1.880 ;
        RECT  12.530 1.540 14.505 1.880 ;
        RECT  14.275 1.540 14.505 3.550 ;
        RECT  13.820 3.320 14.505 3.550 ;
        RECT  13.820 3.320 14.050 4.160 ;
        RECT  13.710 3.820 14.050 4.160 ;
        RECT  1.255 1.585 2.60 1.815 ;
        RECT  4.445 2.870 5.40 3.155 ;
        RECT  4.445 2.925 6.80 3.155 ;
        RECT  2.255 0.630 3.40 0.860 ;
        RECT  10.715 0.630 12.40 0.860 ;
    END
END SDFRRQX1

MACRO SDFRRQX0
    CLASS CORE ;
    FOREIGN SDFRRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.550  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.300 3.010 14.995 3.350 ;
        RECT  14.570 2.860 14.995 3.350 ;
        RECT  14.570 0.630 14.800 3.350 ;
        RECT  14.200 0.630 14.800 0.970 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.830 2.215 9.325 2.720 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.610 2.250 13.105 2.895 ;
        END
    END RN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.300 3.810 14.640 5.280 ;
        RECT  12.285 3.910 12.620 5.280 ;
        RECT  9.510 3.630 9.850 5.280 ;
        RECT  8.310 3.910 8.650 5.280 ;
        RECT  4.830 3.865 5.170 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.400 -0.400 13.740 0.950 ;
        RECT  8.615 -0.400 8.900 1.400 ;
        RECT  4.485 -0.400 4.825 0.655 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  3.500 1.345 5.425 1.575 ;
        RECT  3.505 1.805 5.520 2.090 ;
        RECT  5.235 1.805 5.520 2.180 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.750 1.230 6.655 1.540 ;
        RECT  3.965 2.325 4.950 2.665 ;
        RECT  4.605 2.325 4.950 3.175 ;
        RECT  4.605 2.945 5.980 3.175 ;
        RECT  5.750 1.230 5.980 3.175 ;
        RECT  5.790 3.025 6.500 3.255 ;
        RECT  6.270 3.025 6.500 3.790 ;
        RECT  6.270 3.450 6.610 3.790 ;
        RECT  4.370 3.405 5.615 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.420 3.440 5.650 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.030 3.910 7.370 4.250 ;
        RECT  5.420 4.020 7.370 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  3.960 0.630 4.190 1.115 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  5.290 0.770 7.455 1.000 ;
        RECT  3.960 0.885 5.520 1.115 ;
        RECT  7.115 0.770 7.455 1.570 ;
        RECT  7.875 2.360 8.310 2.700 ;
        RECT  6.210 2.565 7.075 2.795 ;
        RECT  9.590 1.230 9.820 3.330 ;
        RECT  8.080 2.990 10.800 3.330 ;
        RECT  10.455 2.990 10.800 3.395 ;
        RECT  6.845 2.565 7.075 3.680 ;
        RECT  8.080 2.360 8.310 3.680 ;
        RECT  6.845 3.450 8.310 3.680 ;
        RECT  9.130 0.770 10.280 1.000 ;
        RECT  7.815 1.230 8.155 1.870 ;
        RECT  7.815 1.640 9.360 1.870 ;
        RECT  9.130 0.770 9.360 1.870 ;
        RECT  6.210 1.840 8.045 2.110 ;
        RECT  6.210 1.840 7.645 2.180 ;
        RECT  10.050 0.770 10.280 2.425 ;
        RECT  10.050 2.195 10.800 2.425 ;
        RECT  10.460 2.235 11.595 2.535 ;
        RECT  7.415 1.840 7.645 3.220 ;
        RECT  7.415 2.925 7.825 3.220 ;
        RECT  7.415 2.930 7.850 3.220 ;
        RECT  11.255 2.235 11.595 3.440 ;
        RECT  10.510 0.630 12.850 0.860 ;
        RECT  10.510 0.630 10.795 0.970 ;
        RECT  12.510 0.630 12.850 0.970 ;
        RECT  11.485 1.175 12.055 1.515 ;
        RECT  12.805 3.125 13.610 3.465 ;
        RECT  11.825 3.235 13.610 3.465 ;
        RECT  10.805 3.640 11.140 3.970 ;
        RECT  10.805 3.655 11.145 3.970 ;
        RECT  11.825 1.175 12.055 3.970 ;
        RECT  10.805 3.685 12.055 3.970 ;
        RECT  13.840 1.410 14.340 1.750 ;
        RECT  12.450 1.695 14.070 2.020 ;
        RECT  13.840 1.410 14.070 4.175 ;
        RECT  13.195 3.835 14.070 4.175 ;
        RECT  0.980 1.585 2.30 1.960 ;
        RECT  1.445 1.125 2.20 1.355 ;
        RECT  3.505 1.805 4.80 2.090 ;
        RECT  1.995 3.710 3.80 3.940 ;
        RECT  1.980 0.630 3.80 0.860 ;
        RECT  5.290 0.770 6.30 1.000 ;
        RECT  8.080 2.990 9.70 3.330 ;
        RECT  10.510 0.630 11.30 0.860 ;
    END
END SDFRRQX0

MACRO SDFRQX4
    CLASS CORE ;
    FOREIGN SDFRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 1.240 16.830 4.130 ;
        RECT  15.170 2.250 16.830 2.630 ;
        RECT  15.170 0.790 15.510 2.630 ;
        RECT  15.050 2.890 15.400 4.130 ;
        RECT  15.170 0.790 15.400 4.130 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.275 1.640 9.070 2.100 ;
        END
    END C
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.930 -0.400 16.270 0.720 ;
        RECT  14.410 -0.400 14.750 0.710 ;
        RECT  13.005 -0.400 13.345 1.450 ;
        RECT  10.420 -0.400 10.760 1.370 ;
        RECT  8.415 -0.400 8.700 0.950 ;
        RECT  3.485 -0.400 4.935 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 3.470 16.110 5.280 ;
        RECT  14.290 4.160 14.630 5.280 ;
        RECT  12.960 3.530 13.300 5.280 ;
        RECT  10.940 3.965 11.280 5.280 ;
        RECT  8.545 2.910 8.830 5.280 ;
        RECT  4.475 3.965 4.815 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.960 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.400 5.335 1.740 ;
        RECT  3.895 1.400 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.070 1.190 6.395 1.530 ;
        RECT  5.620 1.300 6.395 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  5.620 1.300 5.850 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  5.620 2.935 6.045 3.275 ;
        RECT  4.630 3.045 6.045 3.275 ;
        RECT  6.425 2.980 6.765 3.735 ;
        RECT  2.020 3.505 6.765 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.165 0.730 6.855 0.960 ;
        RECT  2.255 0.940 5.395 1.170 ;
        RECT  6.625 0.730 6.855 1.660 ;
        RECT  6.625 1.320 7.210 1.660 ;
        RECT  8.930 0.775 10.190 1.005 ;
        RECT  7.085 0.735 7.955 1.090 ;
        RECT  7.595 0.735 7.955 1.410 ;
        RECT  8.930 0.775 9.160 1.410 ;
        RECT  7.595 1.180 9.160 1.410 ;
        RECT  9.960 0.775 10.190 1.960 ;
        RECT  9.960 1.730 11.670 1.960 ;
        RECT  11.330 1.730 11.670 2.070 ;
        RECT  7.595 0.735 7.855 2.940 ;
        RECT  6.080 1.840 6.390 2.195 ;
        RECT  6.080 1.965 7.365 2.195 ;
        RECT  9.390 1.240 9.730 2.680 ;
        RECT  9.390 2.340 10.310 2.680 ;
        RECT  12.000 1.540 12.285 2.680 ;
        RECT  8.085 2.450 12.285 2.680 ;
        RECT  9.210 2.450 9.550 2.860 ;
        RECT  7.025 1.965 7.365 3.400 ;
        RECT  8.085 2.450 8.315 3.400 ;
        RECT  7.025 3.170 8.315 3.400 ;
        RECT  9.210 2.450 9.440 3.855 ;
        RECT  10.410 3.505 11.750 3.735 ;
        RECT  9.210 3.625 10.640 3.855 ;
        RECT  11.520 3.650 12.030 3.990 ;
        RECT  11.570 0.970 11.910 1.310 ;
        RECT  11.570 1.080 12.745 1.310 ;
        RECT  13.350 2.355 13.690 2.700 ;
        RECT  12.515 2.470 13.690 2.700 ;
        RECT  12.515 1.080 12.745 3.220 ;
        RECT  9.750 2.990 12.745 3.220 ;
        RECT  11.930 2.990 12.270 3.330 ;
        RECT  9.750 2.990 10.090 3.395 ;
        RECT  13.830 1.070 14.170 1.910 ;
        RECT  12.975 1.680 14.170 1.910 ;
        RECT  12.975 1.680 13.260 2.030 ;
        RECT  13.940 1.070 14.170 3.160 ;
        RECT  13.730 2.930 14.070 3.760 ;
        RECT  1.145 1.585 2.70 1.815 ;
        RECT  2.020 3.505 5.10 3.735 ;
        RECT  2.255 0.940 4.30 1.170 ;
        RECT  8.085 2.450 11.20 2.680 ;
        RECT  9.750 2.990 11.80 3.220 ;
    END
END SDFRQX4

MACRO SDFRQX2
    CLASS CORE ;
    FOREIGN SDFRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.350 1.250 13.735 3.770 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.260 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.680 1.005 2.200 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.130 2.020 8.695 2.630 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.910 -0.400 14.250 0.720 ;
        RECT  12.790 -0.400 13.130 0.720 ;
        RECT  11.385 -0.400 11.730 0.970 ;
        RECT  9.585 -0.400 9.925 0.790 ;
        RECT  7.560 -0.400 7.845 1.330 ;
        RECT  4.100 -0.400 4.440 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.910 4.170 14.250 5.280 ;
        RECT  12.795 4.170 13.135 5.280 ;
        RECT  11.185 3.960 11.525 5.280 ;
        RECT  9.005 3.660 9.345 5.280 ;
        RECT  7.705 3.530 8.045 5.280 ;
        RECT  4.415 4.100 4.755 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.160 2.015 ;
        RECT  4.890 1.785 5.160 2.485 ;
        RECT  3.480 1.400 3.710 3.240 ;
        RECT  3.480 2.900 4.200 3.240 ;
        RECT  5.330 1.205 5.670 1.545 ;
        RECT  3.940 2.245 4.660 2.585 ;
        RECT  4.430 2.245 4.660 2.945 ;
        RECT  4.430 2.715 5.620 2.945 ;
        RECT  5.390 1.205 5.620 3.385 ;
        RECT  5.390 3.045 5.985 3.385 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  4.690 0.745 6.470 0.975 ;
        RECT  1.770 0.940 4.920 1.170 ;
        RECT  6.130 0.745 6.470 1.595 ;
        RECT  6.405 3.530 6.745 3.870 ;
        RECT  2.120 3.640 6.745 3.870 ;
        RECT  2.120 3.640 2.410 4.020 ;
        RECT  8.075 0.680 9.355 0.910 ;
        RECT  6.785 0.630 7.125 0.965 ;
        RECT  9.125 0.680 9.355 1.250 ;
        RECT  9.125 1.020 9.615 1.250 ;
        RECT  9.385 1.020 9.615 1.920 ;
        RECT  8.075 0.680 8.305 1.790 ;
        RECT  6.895 1.560 8.305 1.790 ;
        RECT  9.385 1.690 10.550 1.920 ;
        RECT  10.210 1.690 10.550 2.100 ;
        RECT  6.895 0.630 7.125 2.165 ;
        RECT  6.520 1.825 7.285 2.165 ;
        RECT  6.945 1.560 7.285 2.825 ;
        RECT  8.535 1.140 8.895 1.480 ;
        RECT  8.665 1.480 9.155 1.710 ;
        RECT  5.850 1.900 6.190 2.625 ;
        RECT  5.850 2.395 6.445 2.625 ;
        RECT  9.675 2.360 11.060 2.700 ;
        RECT  8.925 2.470 11.060 2.700 ;
        RECT  7.515 2.020 7.800 3.300 ;
        RECT  6.215 2.395 6.445 3.300 ;
        RECT  7.515 2.960 9.155 3.300 ;
        RECT  8.925 1.480 9.155 3.300 ;
        RECT  6.215 3.055 9.155 3.300 ;
        RECT  10.560 0.630 10.900 0.970 ;
        RECT  10.670 0.630 10.900 1.460 ;
        RECT  10.670 1.230 11.520 1.460 ;
        RECT  11.290 1.230 11.520 3.160 ;
        RECT  12.370 2.340 12.655 3.160 ;
        RECT  10.155 2.930 12.655 3.160 ;
        RECT  10.155 2.930 10.495 3.825 ;
        RECT  12.090 0.680 12.430 2.105 ;
        RECT  11.750 1.875 13.115 2.105 ;
        RECT  11.750 1.875 12.040 2.650 ;
        RECT  12.885 1.875 13.115 3.730 ;
        RECT  12.030 3.390 13.115 3.730 ;
        RECT  1.770 0.940 3.60 1.170 ;
        RECT  2.120 3.640 5.60 3.870 ;
        RECT  8.925 2.470 10.90 2.700 ;
        RECT  6.215 3.055 8.80 3.300 ;
        RECT  10.155 2.930 11.20 3.160 ;
    END
END SDFRQX2

MACRO SDFRQX1
    CLASS CORE ;
    FOREIGN SDFRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.420 2.250 14.375 2.630 ;
        RECT  13.160 3.780 13.650 4.120 ;
        RECT  13.420 0.700 13.650 4.120 ;
        RECT  13.160 0.700 13.650 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 3.990 2.030 4.250 ;
        RECT  1.610 3.980 2.000 4.250 ;
        RECT  1.610 3.470 1.840 4.250 ;
        RECT  1.410 3.470 1.840 3.815 ;
        RECT  1.385 3.470 1.840 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.880 2.800 3.655 3.240 ;
        RECT  2.880 2.045 3.110 3.240 ;
        RECT  0.575 2.045 3.110 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 1.640 8.885 2.035 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.880 -0.400 14.220 1.040 ;
        RECT  12.000 -0.400 12.340 1.030 ;
        RECT  10.145 -0.400 10.485 1.030 ;
        RECT  8.085 -0.400 8.425 0.950 ;
        RECT  4.725 -0.400 5.065 0.655 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  2.825 1.090 3.825 1.320 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.880 3.330 14.220 5.280 ;
        RECT  12.365 4.040 12.705 5.280 ;
        RECT  9.480 3.500 9.820 5.280 ;
        RECT  8.180 3.620 8.520 5.280 ;
        RECT  4.905 3.845 5.230 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.630 1.815 ;
        RECT  3.290 1.555 3.630 1.895 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  3.900 1.755 4.240 2.110 ;
        RECT  3.900 1.880 5.275 2.110 ;
        RECT  4.935 1.880 5.275 2.220 ;
        RECT  3.900 1.755 4.215 3.425 ;
        RECT  5.885 1.200 6.225 1.540 ;
        RECT  4.445 2.565 4.775 3.155 ;
        RECT  5.680 1.310 5.920 3.155 ;
        RECT  4.445 2.925 6.460 3.155 ;
        RECT  6.120 2.925 6.460 3.460 ;
        RECT  2.255 0.630 4.495 0.860 ;
        RECT  4.265 0.630 4.495 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.295 0.740 7.025 0.970 ;
        RECT  4.265 0.885 5.525 1.115 ;
        RECT  6.685 0.740 7.025 1.685 ;
        RECT  2.070 3.420 2.410 3.760 ;
        RECT  4.445 3.385 5.710 3.615 ;
        RECT  5.480 3.385 5.710 3.930 ;
        RECT  2.070 3.530 3.580 3.760 ;
        RECT  4.445 3.385 4.675 3.885 ;
        RECT  3.365 3.655 4.675 3.885 ;
        RECT  6.880 3.620 7.220 3.930 ;
        RECT  5.480 3.700 7.220 3.930 ;
        RECT  9.115 1.095 9.455 1.460 ;
        RECT  6.165 2.165 6.505 2.675 ;
        RECT  7.745 2.105 8.095 2.460 ;
        RECT  6.165 2.445 7.010 2.675 ;
        RECT  9.115 1.095 9.345 3.230 ;
        RECT  8.940 2.710 9.345 3.230 ;
        RECT  6.780 2.445 7.010 3.390 ;
        RECT  7.990 2.245 8.220 3.390 ;
        RECT  8.940 2.890 10.730 3.230 ;
        RECT  6.780 3.160 9.170 3.390 ;
        RECT  8.655 0.630 9.915 0.860 ;
        RECT  7.285 0.645 7.625 1.410 ;
        RECT  8.655 0.630 8.885 1.410 ;
        RECT  7.285 1.180 8.885 1.410 ;
        RECT  6.965 1.915 7.515 2.205 ;
        RECT  9.685 0.630 9.915 2.450 ;
        RECT  9.685 2.220 10.465 2.450 ;
        RECT  10.125 2.330 11.210 2.560 ;
        RECT  7.285 0.645 7.515 2.930 ;
        RECT  7.285 2.690 7.760 2.930 ;
        RECT  10.980 2.330 11.210 3.320 ;
        RECT  10.980 2.980 11.405 3.320 ;
        RECT  10.995 0.710 11.670 1.070 ;
        RECT  11.440 2.430 11.885 2.660 ;
        RECT  11.440 0.710 11.670 2.660 ;
        RECT  11.650 2.660 12.520 3.000 ;
        RECT  10.630 3.545 10.930 3.840 ;
        RECT  10.740 3.550 10.970 4.215 ;
        RECT  11.650 2.430 11.880 4.215 ;
        RECT  10.740 3.985 11.880 4.215 ;
        RECT  11.900 1.615 13.140 1.955 ;
        RECT  11.900 1.615 12.185 2.135 ;
        RECT  12.910 1.615 13.140 3.470 ;
        RECT  12.460 3.240 13.140 3.470 ;
        RECT  12.460 3.240 12.800 3.580 ;
        RECT  1.255 1.585 2.80 1.815 ;
        RECT  4.445 2.925 5.30 3.155 ;
        RECT  2.255 0.630 3.70 0.860 ;
        RECT  6.780 3.160 8.30 3.390 ;
    END
END SDFRQX1

MACRO SDFRQX0
    CLASS CORE ;
    FOREIGN SDFRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 1.640 13.105 2.020 ;
        RECT  12.620 3.430 12.960 3.770 ;
        RECT  12.725 1.640 12.960 3.770 ;
        RECT  12.725 0.630 12.955 3.770 ;
        RECT  12.045 0.630 12.955 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.215 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.215 3.320 ;
        RECT  2.190 2.860 3.215 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.625 2.185 8.120 2.675 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  12.020 4.165 12.360 5.280 ;
        RECT  10.755 3.910 11.040 5.280 ;
        RECT  7.650 3.650 8.460 5.280 ;
        RECT  3.200 4.170 4.495 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  9.270 -0.400 9.555 0.710 ;
        RECT  9.250 -0.400 9.555 0.675 ;
        RECT  7.375 -0.400 7.660 0.970 ;
        RECT  3.970 -0.400 4.310 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.215 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.445 1.805 4.770 2.035 ;
        RECT  3.445 1.805 3.875 2.095 ;
        RECT  3.445 1.805 3.835 2.105 ;
        RECT  4.485 1.805 4.770 2.205 ;
        RECT  3.445 1.805 3.675 3.425 ;
        RECT  3.445 3.085 4.195 3.425 ;
        RECT  5.000 1.230 5.800 1.540 ;
        RECT  3.905 2.325 4.190 2.665 ;
        RECT  3.905 2.435 5.230 2.665 ;
        RECT  5.000 1.230 5.230 3.480 ;
        RECT  4.995 2.435 5.230 3.480 ;
        RECT  4.995 3.250 5.725 3.480 ;
        RECT  5.385 3.250 5.725 3.790 ;
        RECT  1.995 3.710 5.050 3.940 ;
        RECT  4.820 3.710 5.050 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.145 3.925 6.485 4.250 ;
        RECT  4.820 4.020 6.485 4.250 ;
        RECT  4.540 0.630 6.500 0.920 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  4.540 0.630 4.770 1.355 ;
        RECT  1.980 1.125 4.770 1.355 ;
        RECT  5.460 2.440 5.800 2.780 ;
        RECT  7.045 2.355 7.395 2.695 ;
        RECT  5.460 2.530 6.190 2.780 ;
        RECT  8.350 2.605 9.410 2.945 ;
        RECT  8.350 1.230 8.580 3.245 ;
        RECT  7.165 2.905 8.580 3.245 ;
        RECT  5.960 2.530 6.190 3.695 ;
        RECT  7.165 2.355 7.395 3.695 ;
        RECT  5.960 3.465 7.395 3.695 ;
        RECT  7.890 0.770 9.040 1.000 ;
        RECT  7.890 0.770 8.120 1.480 ;
        RECT  6.865 1.250 8.120 1.480 ;
        RECT  8.810 0.770 9.040 2.165 ;
        RECT  6.865 1.250 7.205 2.110 ;
        RECT  5.460 1.770 7.205 2.110 ;
        RECT  8.810 1.935 9.580 2.165 ;
        RECT  9.240 2.045 10.065 2.275 ;
        RECT  6.585 1.770 6.815 3.230 ;
        RECT  6.585 2.895 6.930 3.230 ;
        RECT  6.585 2.900 6.935 3.230 ;
        RECT  9.725 2.045 10.065 3.400 ;
        RECT  10.125 1.110 10.525 1.450 ;
        RECT  11.390 2.370 11.730 2.710 ;
        RECT  10.295 2.480 11.730 2.710 ;
        RECT  10.295 1.110 10.525 3.970 ;
        RECT  9.350 3.650 10.525 3.970 ;
        RECT  12.045 1.350 12.385 1.900 ;
        RECT  11.085 1.700 12.190 2.040 ;
        RECT  11.960 1.700 12.190 3.565 ;
        RECT  11.220 3.225 12.190 3.565 ;
        RECT  0.980 1.585 2.70 1.960 ;
        RECT  1.995 3.710 4.90 3.940 ;
        RECT  1.980 1.125 3.70 1.355 ;
    END
END SDFRQX0

MACRO SDFFX4
    CLASS CORE ;
    FOREIGN SDFFX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.290  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.010 1.130 19.350 4.100 ;
        RECT  17.680 2.250 19.350 2.630 ;
        RECT  17.680 2.250 18.030 3.770 ;
        RECT  17.680 1.130 17.910 3.770 ;
        RECT  17.570 1.130 17.910 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.980 2.885 17.410 3.115 ;
        RECT  17.180 1.700 17.410 3.115 ;
        RECT  14.690 1.700 17.410 1.930 ;
        RECT  16.420 2.885 16.760 4.130 ;
        RECT  16.130 1.130 16.470 1.930 ;
        RECT  14.980 2.885 16.760 3.240 ;
        RECT  14.980 2.860 15.625 3.240 ;
        RECT  14.980 2.860 15.320 4.130 ;
        RECT  14.690 1.130 15.030 1.930 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.275 1.640 9.070 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.290 -0.400 18.630 1.470 ;
        RECT  16.850 -0.400 17.190 1.470 ;
        RECT  15.410 -0.400 15.750 1.470 ;
        RECT  13.095 -0.400 13.435 1.450 ;
        RECT  10.420 -0.400 10.760 1.370 ;
        RECT  8.415 -0.400 8.700 0.950 ;
        RECT  3.485 -0.400 4.935 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.250 4.170 18.590 5.280 ;
        RECT  17.130 4.170 17.470 5.280 ;
        RECT  15.700 3.470 16.040 5.280 ;
        RECT  14.220 4.160 14.560 5.280 ;
        RECT  12.960 3.770 13.300 5.280 ;
        RECT  10.940 4.225 11.280 5.280 ;
        RECT  8.545 2.910 8.830 5.280 ;
        RECT  4.475 3.965 4.815 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.960 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.400 5.335 1.740 ;
        RECT  3.895 1.400 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.070 1.190 6.395 1.530 ;
        RECT  5.620 1.300 6.395 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  5.620 1.300 5.850 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  5.620 2.935 6.045 3.275 ;
        RECT  4.630 3.045 6.045 3.275 ;
        RECT  6.425 2.980 6.765 3.735 ;
        RECT  2.020 3.505 6.765 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  5.165 0.630 6.855 0.860 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.165 0.630 5.395 1.170 ;
        RECT  2.255 0.940 5.395 1.170 ;
        RECT  6.625 0.630 6.855 1.660 ;
        RECT  6.625 1.320 7.210 1.660 ;
        RECT  8.930 0.775 10.190 1.005 ;
        RECT  7.595 0.735 7.955 1.410 ;
        RECT  8.930 0.775 9.160 1.410 ;
        RECT  7.595 1.180 9.160 1.410 ;
        RECT  12.000 1.440 12.340 1.780 ;
        RECT  6.080 1.840 6.390 2.195 ;
        RECT  6.080 1.965 7.855 2.195 ;
        RECT  9.960 0.775 10.190 2.940 ;
        RECT  7.595 0.735 7.855 2.940 ;
        RECT  12.000 1.440 12.230 2.940 ;
        RECT  9.960 2.600 12.230 2.940 ;
        RECT  9.390 1.240 9.730 2.680 ;
        RECT  8.085 2.450 9.730 2.680 ;
        RECT  7.025 2.545 7.365 3.400 ;
        RECT  8.085 2.450 8.315 3.400 ;
        RECT  7.025 3.170 8.315 3.400 ;
        RECT  9.210 2.450 9.520 4.115 ;
        RECT  10.410 3.765 11.750 3.995 ;
        RECT  9.210 3.885 10.640 4.115 ;
        RECT  11.520 3.945 12.550 4.175 ;
        RECT  11.570 0.870 11.910 1.210 ;
        RECT  11.570 0.980 12.800 1.210 ;
        RECT  13.460 2.355 13.800 2.700 ;
        RECT  12.570 2.470 13.800 2.700 ;
        RECT  12.570 0.980 12.800 3.480 ;
        RECT  9.750 3.250 12.800 3.480 ;
        RECT  11.930 3.250 12.270 3.590 ;
        RECT  9.750 3.250 10.090 3.655 ;
        RECT  13.940 1.070 14.280 1.910 ;
        RECT  13.030 1.680 14.280 1.910 ;
        RECT  13.030 1.680 13.370 2.030 ;
        RECT  14.050 2.310 16.950 2.540 ;
        RECT  16.610 2.310 16.950 2.650 ;
        RECT  14.050 1.070 14.280 3.160 ;
        RECT  13.660 2.930 14.280 3.160 ;
        RECT  13.660 2.930 14.000 3.760 ;
        RECT  1.145 1.585 2.80 1.815 ;
        RECT  2.020 3.505 5.30 3.735 ;
        RECT  2.255 0.940 4.20 1.170 ;
        RECT  9.960 2.600 11.80 2.940 ;
        RECT  9.750 3.250 11.60 3.480 ;
        RECT  14.050 2.310 15.40 2.540 ;
    END
END SDFFX4

MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.350 3.270 14.365 3.500 ;
        RECT  14.135 1.250 14.365 3.500 ;
        RECT  13.985 2.860 14.365 3.500 ;
        RECT  13.350 1.250 14.365 1.590 ;
        RECT  13.350 3.270 13.690 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.260 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.620 1.890 4.250 ;
        RECT  0.755 3.620 1.890 3.850 ;
        RECT  0.755 3.470 1.135 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.720 1.005 2.200 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 1.240 15.010 3.550 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.130 2.020 8.695 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.230 -0.400 15.570 0.720 ;
        RECT  14.110 -0.400 14.450 0.720 ;
        RECT  12.790 -0.400 13.130 0.720 ;
        RECT  11.385 -0.400 11.730 0.970 ;
        RECT  9.585 -0.400 9.925 0.790 ;
        RECT  7.560 -0.400 7.845 1.330 ;
        RECT  4.100 -0.400 4.440 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.230 3.950 15.570 5.280 ;
        RECT  14.110 3.950 14.450 5.280 ;
        RECT  12.590 4.125 12.930 5.280 ;
        RECT  11.185 3.990 11.525 5.280 ;
        RECT  9.005 3.690 9.345 5.280 ;
        RECT  7.705 3.530 8.045 5.280 ;
        RECT  4.415 4.100 4.755 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.160 2.015 ;
        RECT  4.890 1.785 5.160 2.485 ;
        RECT  3.480 1.400 3.710 3.240 ;
        RECT  3.480 2.900 4.200 3.240 ;
        RECT  5.330 1.205 5.670 1.545 ;
        RECT  3.940 2.245 4.660 2.585 ;
        RECT  4.430 2.245 4.660 2.945 ;
        RECT  4.430 2.715 5.620 2.945 ;
        RECT  5.390 1.205 5.620 3.385 ;
        RECT  5.390 3.045 5.985 3.385 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  4.690 0.745 6.470 0.975 ;
        RECT  1.770 0.940 4.920 1.170 ;
        RECT  6.130 0.745 6.470 1.595 ;
        RECT  6.405 3.220 6.745 3.870 ;
        RECT  2.120 3.640 6.745 3.870 ;
        RECT  2.120 3.640 2.410 4.020 ;
        RECT  8.075 0.680 9.355 0.910 ;
        RECT  6.785 0.630 7.125 0.965 ;
        RECT  9.125 0.680 9.355 1.250 ;
        RECT  9.125 1.020 9.615 1.250 ;
        RECT  6.895 0.630 7.125 1.790 ;
        RECT  8.075 0.680 8.305 1.790 ;
        RECT  6.895 1.560 8.305 1.790 ;
        RECT  9.385 1.020 9.615 2.460 ;
        RECT  5.850 1.900 6.190 2.625 ;
        RECT  9.385 2.120 9.755 2.460 ;
        RECT  5.850 2.395 7.285 2.625 ;
        RECT  6.945 1.560 7.285 2.880 ;
        RECT  8.535 1.140 8.895 1.710 ;
        RECT  8.535 1.480 9.155 1.710 ;
        RECT  10.210 1.720 10.550 3.255 ;
        RECT  7.515 2.020 7.800 3.255 ;
        RECT  8.925 1.480 9.155 3.255 ;
        RECT  7.515 2.915 9.155 3.255 ;
        RECT  10.210 2.820 10.685 3.255 ;
        RECT  7.515 3.025 10.685 3.255 ;
        RECT  10.560 0.630 10.900 0.970 ;
        RECT  10.670 0.630 10.900 1.460 ;
        RECT  10.670 1.230 11.520 1.460 ;
        RECT  12.370 2.750 12.655 3.160 ;
        RECT  11.290 2.930 12.655 3.160 ;
        RECT  11.290 1.230 11.520 3.715 ;
        RECT  10.155 3.485 11.520 3.715 ;
        RECT  10.155 3.485 10.495 3.825 ;
        RECT  12.090 0.680 12.430 2.520 ;
        RECT  11.750 2.290 13.380 2.520 ;
        RECT  11.750 2.290 12.040 2.650 ;
        RECT  12.885 2.290 13.380 2.650 ;
        RECT  12.885 2.290 13.115 3.720 ;
        RECT  12.030 3.390 13.115 3.720 ;
        RECT  1.770 0.940 3.90 1.170 ;
        RECT  2.120 3.640 5.40 3.870 ;
        RECT  7.515 3.025 9.60 3.255 ;
    END
END SDFFX2

MACRO SDFFX1
    CLASS CORE ;
    FOREIGN SDFFX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.605 0.940 14.995 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 1.640 14.375 2.020 ;
        RECT  13.420 2.870 14.220 3.100 ;
        RECT  13.985 1.640 14.220 3.100 ;
        RECT  13.985 1.260 14.215 3.100 ;
        RECT  13.420 1.260 14.215 1.490 ;
        RECT  13.160 3.780 13.650 4.120 ;
        RECT  13.420 2.870 13.650 4.120 ;
        RECT  13.420 0.700 13.650 1.490 ;
        RECT  13.160 0.700 13.650 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 3.990 2.030 4.250 ;
        RECT  1.610 3.980 2.000 4.250 ;
        RECT  1.610 3.470 1.840 4.250 ;
        RECT  1.410 3.470 1.840 3.815 ;
        RECT  1.385 3.470 1.840 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.880 2.800 3.655 3.240 ;
        RECT  2.880 2.045 3.110 3.240 ;
        RECT  0.575 2.045 3.110 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 1.640 8.885 2.035 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.880 -0.400 14.220 1.030 ;
        RECT  12.000 -0.400 12.340 1.020 ;
        RECT  10.145 -0.400 10.485 0.710 ;
        RECT  8.085 -0.400 8.425 0.950 ;
        RECT  4.725 -0.400 5.065 0.655 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  2.825 1.090 3.825 1.320 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  13.880 3.330 14.220 5.280 ;
        RECT  12.365 4.040 12.705 5.280 ;
        RECT  9.480 3.620 9.820 5.280 ;
        RECT  8.180 2.725 8.520 5.280 ;
        RECT  4.905 3.845 5.230 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.630 1.815 ;
        RECT  3.290 1.555 3.630 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  3.900 1.755 4.240 2.110 ;
        RECT  3.900 1.880 5.275 2.110 ;
        RECT  4.935 1.880 5.275 2.220 ;
        RECT  3.900 1.755 4.215 3.425 ;
        RECT  5.885 1.200 6.225 1.540 ;
        RECT  4.445 2.565 4.775 3.155 ;
        RECT  5.680 1.310 5.920 3.155 ;
        RECT  4.445 2.925 6.460 3.155 ;
        RECT  6.120 2.925 6.460 3.460 ;
        RECT  2.255 0.630 4.495 0.860 ;
        RECT  4.265 0.630 4.495 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.295 0.740 7.025 0.970 ;
        RECT  4.265 0.885 5.525 1.115 ;
        RECT  6.685 0.740 7.025 1.685 ;
        RECT  2.070 3.420 2.410 3.760 ;
        RECT  4.445 3.385 5.710 3.615 ;
        RECT  5.480 3.385 5.710 3.930 ;
        RECT  2.070 3.530 3.580 3.760 ;
        RECT  4.445 3.385 4.675 3.885 ;
        RECT  3.365 3.655 4.675 3.885 ;
        RECT  6.880 3.320 7.220 3.930 ;
        RECT  5.480 3.700 7.220 3.930 ;
        RECT  8.655 0.630 9.915 0.860 ;
        RECT  7.285 0.645 7.625 1.410 ;
        RECT  8.655 0.630 8.885 1.410 ;
        RECT  7.285 1.180 8.885 1.410 ;
        RECT  6.165 2.165 6.505 2.505 ;
        RECT  6.165 2.275 7.515 2.505 ;
        RECT  9.685 0.630 9.915 2.885 ;
        RECT  7.285 0.645 7.515 2.975 ;
        RECT  9.685 2.575 10.730 2.885 ;
        RECT  7.285 2.690 7.760 2.975 ;
        RECT  9.115 1.095 9.455 1.460 ;
        RECT  10.185 1.900 10.525 2.240 ;
        RECT  10.185 2.010 11.210 2.240 ;
        RECT  7.745 2.245 8.220 2.460 ;
        RECT  7.745 2.105 8.095 2.460 ;
        RECT  7.990 2.265 9.345 2.495 ;
        RECT  10.980 2.010 11.210 3.345 ;
        RECT  9.115 1.095 9.345 3.345 ;
        RECT  8.940 2.265 9.345 3.345 ;
        RECT  10.980 2.980 11.405 3.345 ;
        RECT  8.940 3.115 11.405 3.345 ;
        RECT  10.995 0.710 11.670 1.070 ;
        RECT  11.440 2.430 11.885 2.660 ;
        RECT  11.440 0.710 11.670 2.660 ;
        RECT  11.650 2.660 12.520 3.000 ;
        RECT  11.650 2.430 11.880 3.960 ;
        RECT  10.630 3.615 11.880 3.960 ;
        RECT  11.900 1.615 13.195 1.955 ;
        RECT  12.960 1.615 13.195 2.475 ;
        RECT  11.900 1.615 12.185 2.135 ;
        RECT  12.960 2.135 13.355 2.475 ;
        RECT  12.960 1.615 13.190 3.470 ;
        RECT  12.460 3.240 13.190 3.470 ;
        RECT  12.460 3.240 12.800 3.580 ;
        RECT  1.255 1.585 2.50 1.815 ;
        RECT  4.445 2.925 5.30 3.155 ;
        RECT  2.255 0.630 3.40 0.860 ;
        RECT  8.940 3.115 10.60 3.345 ;
    END
END SDFFX1

MACRO SDFFX0
    CLASS CORE ;
    FOREIGN SDFFX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.220 2.860 13.735 3.240 ;
        RECT  13.220 2.640 13.640 3.240 ;
        RECT  13.410 1.170 13.640 3.240 ;
        RECT  13.300 1.170 13.640 1.510 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.602  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 1.640 13.105 2.020 ;
        RECT  12.330 2.710 12.955 3.050 ;
        RECT  12.725 0.630 12.955 3.050 ;
        RECT  12.045 0.630 12.955 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.215 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.215 3.320 ;
        RECT  2.190 2.860 3.215 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.625 2.185 8.120 2.675 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  13.220 3.470 13.560 5.280 ;
        RECT  11.730 4.165 12.070 5.280 ;
        RECT  10.755 4.040 11.040 5.280 ;
        RECT  8.120 3.630 8.460 5.280 ;
        RECT  7.395 3.850 7.735 5.280 ;
        RECT  3.200 4.170 4.495 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.300 -0.400 13.640 0.710 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  9.270 -0.400 9.555 0.710 ;
        RECT  9.250 -0.400 9.555 0.675 ;
        RECT  7.375 -0.400 7.660 0.970 ;
        RECT  3.970 -0.400 4.310 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.215 1.815 ;
        RECT  2.930 1.585 3.215 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.445 1.805 4.770 2.035 ;
        RECT  3.445 1.805 3.875 2.105 ;
        RECT  4.485 1.805 4.770 2.205 ;
        RECT  3.445 1.805 3.675 3.425 ;
        RECT  3.445 3.085 4.195 3.425 ;
        RECT  5.000 1.230 5.800 1.540 ;
        RECT  3.905 2.380 4.190 2.720 ;
        RECT  3.905 2.490 5.230 2.720 ;
        RECT  5.000 1.230 5.230 3.480 ;
        RECT  4.995 2.490 5.230 3.480 ;
        RECT  4.995 3.250 5.725 3.480 ;
        RECT  5.385 3.250 5.725 3.790 ;
        RECT  1.995 3.710 5.050 3.940 ;
        RECT  4.820 3.710 5.050 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.145 3.510 6.485 4.250 ;
        RECT  4.820 4.020 6.485 4.250 ;
        RECT  4.540 0.630 6.500 0.860 ;
        RECT  6.160 0.630 6.500 0.970 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  4.540 0.630 4.770 1.355 ;
        RECT  1.980 1.125 4.770 1.355 ;
        RECT  5.460 1.825 6.855 2.165 ;
        RECT  7.890 0.770 9.040 1.000 ;
        RECT  7.890 0.770 8.120 1.480 ;
        RECT  6.865 1.250 8.120 1.480 ;
        RECT  6.865 1.250 7.395 1.590 ;
        RECT  6.705 2.395 7.395 2.625 ;
        RECT  8.810 0.770 9.040 2.885 ;
        RECT  7.165 1.250 7.395 2.625 ;
        RECT  5.845 2.525 6.935 2.865 ;
        RECT  8.810 2.600 9.410 2.885 ;
        RECT  6.585 2.525 6.935 3.155 ;
        RECT  9.295 1.930 9.635 2.270 ;
        RECT  9.295 2.040 9.955 2.270 ;
        RECT  9.725 2.040 9.955 3.400 ;
        RECT  8.350 1.230 8.580 3.345 ;
        RECT  7.995 2.905 8.580 3.345 ;
        RECT  7.165 3.115 10.065 3.345 ;
        RECT  0.980 1.585 2.50 1.815 ;
        RECT  1.995 3.710 4.20 3.940 ;
        RECT  1.980 1.125 3.60 1.355 ;
        RECT  7.165 3.115 9.40 3.345 ;
        RECT  9.725 3.110 10.065 3.400 ;
        RECT  7.165 3.115 7.395 3.620 ;
        RECT  6.875 3.390 7.395 3.620 ;
        RECT  10.125 1.110 10.525 1.450 ;
        RECT  11.300 2.370 11.640 2.710 ;
        RECT  10.295 2.480 11.640 2.710 ;
        RECT  10.295 1.110 10.525 3.970 ;
        RECT  9.350 3.630 10.525 3.970 ;
        RECT  12.045 1.350 12.385 2.320 ;
        RECT  11.085 1.700 12.385 2.040 ;
        RECT  11.870 1.980 12.495 2.320 ;
        RECT  11.130 3.055 11.470 3.455 ;
        RECT  11.870 1.700 12.100 3.455 ;
        RECT  11.130 3.225 12.100 3.455 ;
    END
END SDFFX0

MACRO SDFFSX4
    CLASS CORE ;
    FOREIGN SDFFSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.085  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 1.130 19.980 3.060 ;
        RECT  18.360 2.250 19.980 2.630 ;
        RECT  18.360 2.250 18.715 3.060 ;
        RECT  18.360 1.130 18.590 3.060 ;
        RECT  18.200 1.130 18.590 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.090  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.635 2.880 18.065 3.110 ;
        RECT  17.835 1.700 18.065 3.110 ;
        RECT  15.535 1.700 18.065 1.930 ;
        RECT  15.635 2.880 17.415 3.240 ;
        RECT  16.760 1.130 17.100 1.930 ;
        RECT  15.635 2.860 16.255 3.240 ;
        RECT  15.635 2.860 15.975 4.100 ;
        RECT  15.535 0.700 15.765 1.930 ;
        RECT  15.280 0.700 15.765 1.040 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.760 1.640 14.365 2.070 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 1.640 8.920 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.470 ;
        RECT  17.480 -0.400 17.820 1.470 ;
        RECT  16.040 -0.400 16.380 1.470 ;
        RECT  13.480 -0.400 13.820 0.840 ;
        RECT  10.715 -0.400 11.000 1.370 ;
        RECT  8.820 -0.400 9.105 0.950 ;
        RECT  3.400 -0.400 5.150 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  19.000 3.295 19.340 5.280 ;
        RECT  17.625 3.555 17.965 5.280 ;
        RECT  16.355 3.470 16.695 5.280 ;
        RECT  14.875 4.140 15.215 5.280 ;
        RECT  13.590 2.890 13.930 5.280 ;
        RECT  11.370 3.965 11.710 5.280 ;
        RECT  8.975 2.910 9.260 5.280 ;
        RECT  4.795 3.965 5.135 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.585 5.740 1.875 ;
        RECT  5.400 1.585 5.740 2.265 ;
        RECT  3.895 1.585 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.025 1.190 6.800 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  6.025 1.190 6.255 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  6.025 2.935 6.450 3.275 ;
        RECT  4.630 3.045 6.450 3.275 ;
        RECT  6.830 2.980 7.165 3.735 ;
        RECT  2.020 3.505 7.165 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.380 0.730 7.260 0.960 ;
        RECT  2.255 0.940 5.610 1.170 ;
        RECT  7.030 0.730 7.260 1.660 ;
        RECT  7.030 1.320 7.615 1.660 ;
        RECT  9.335 0.775 10.485 1.005 ;
        RECT  7.490 0.735 8.360 1.090 ;
        RECT  7.855 0.735 8.360 1.410 ;
        RECT  7.855 1.180 9.565 1.410 ;
        RECT  10.255 0.775 10.485 1.960 ;
        RECT  10.255 1.730 11.910 1.960 ;
        RECT  11.570 1.730 11.910 2.070 ;
        RECT  9.335 0.775 9.565 2.100 ;
        RECT  9.210 1.760 9.565 2.100 ;
        RECT  7.855 0.735 8.085 2.940 ;
        RECT  7.855 2.600 8.285 2.940 ;
        RECT  6.485 1.840 6.795 2.195 ;
        RECT  6.485 1.965 7.625 2.195 ;
        RECT  9.795 1.240 10.025 2.680 ;
        RECT  9.795 2.340 10.740 2.680 ;
        RECT  12.240 1.540 12.525 2.680 ;
        RECT  8.515 2.450 12.525 2.680 ;
        RECT  9.640 2.450 9.980 2.860 ;
        RECT  7.395 1.965 7.625 3.400 ;
        RECT  8.515 2.450 8.745 3.400 ;
        RECT  7.395 3.170 8.745 3.400 ;
        RECT  9.640 2.450 9.870 3.855 ;
        RECT  10.840 3.505 12.180 3.735 ;
        RECT  11.950 3.505 12.180 4.100 ;
        RECT  9.640 3.625 11.070 3.855 ;
        RECT  11.950 3.760 12.460 4.100 ;
        RECT  11.810 0.970 12.150 1.310 ;
        RECT  11.810 1.080 12.985 1.310 ;
        RECT  14.505 2.320 14.845 2.660 ;
        RECT  12.755 2.430 14.845 2.660 ;
        RECT  12.755 1.080 12.985 3.220 ;
        RECT  10.180 2.990 12.985 3.220 ;
        RECT  12.360 2.990 12.700 3.330 ;
        RECT  10.180 2.990 10.520 3.395 ;
        RECT  13.215 1.180 15.050 1.410 ;
        RECT  14.710 1.180 15.050 1.700 ;
        RECT  13.215 1.180 13.500 1.530 ;
        RECT  14.710 1.470 15.305 1.700 ;
        RECT  15.075 2.310 17.605 2.540 ;
        RECT  17.265 2.310 17.605 2.650 ;
        RECT  15.075 1.470 15.305 3.120 ;
        RECT  14.315 2.890 15.305 3.120 ;
        RECT  14.315 2.890 14.655 3.730 ;
        RECT  1.145 1.585 2.80 1.815 ;
        RECT  2.020 3.505 6.80 3.735 ;
        RECT  2.255 0.940 4.70 1.170 ;
        RECT  8.515 2.450 11.00 2.680 ;
        RECT  12.755 2.430 13.60 2.660 ;
        RECT  10.180 2.990 11.50 3.220 ;
        RECT  15.075 2.310 16.60 2.540 ;
    END
END SDFFSX4

MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.765 0.830 14.995 3.240 ;
        RECT  14.450 2.860 14.790 4.180 ;
        RECT  14.610 0.830 14.995 1.170 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.720 1.005 2.200 ;
        END
    END SE
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.585 2.050 13.105 2.630 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.875 1.240 16.270 2.020 ;
        RECT  15.770 2.640 16.110 3.550 ;
        RECT  15.875 1.240 16.110 3.550 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.645 1.640 8.115 2.160 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 0.720 ;
        RECT  15.370 -0.400 15.710 0.720 ;
        RECT  13.850 -0.400 14.190 0.970 ;
        RECT  12.300 -0.400 12.645 1.090 ;
        RECT  9.975 -0.400 10.315 0.710 ;
        RECT  8.015 -0.400 8.300 0.950 ;
        RECT  4.530 -0.400 4.870 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.490 2.640 16.830 5.280 ;
        RECT  15.210 3.950 15.550 5.280 ;
        RECT  13.690 4.170 14.030 5.280 ;
        RECT  11.710 3.385 12.750 5.280 ;
        RECT  9.330 3.480 9.670 5.280 ;
        RECT  8.030 3.515 8.370 5.280 ;
        RECT  4.715 3.900 5.055 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.330 2.015 ;
        RECT  4.990 1.785 5.330 2.470 ;
        RECT  3.480 1.400 3.710 3.270 ;
        RECT  3.480 2.930 4.250 3.265 ;
        RECT  3.480 2.930 4.240 3.270 ;
        RECT  5.580 1.190 6.100 1.530 ;
        RECT  3.940 2.245 4.715 2.585 ;
        RECT  4.485 2.245 4.715 2.930 ;
        RECT  5.580 1.190 5.810 3.210 ;
        RECT  4.485 2.700 5.810 2.930 ;
        RECT  5.580 2.870 6.285 3.210 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  5.120 0.730 6.900 0.960 ;
        RECT  1.770 0.940 5.350 1.170 ;
        RECT  6.560 0.730 6.900 1.595 ;
        RECT  4.400 3.440 5.525 3.670 ;
        RECT  2.120 3.500 4.560 3.730 ;
        RECT  5.295 3.515 7.045 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  8.530 0.800 9.735 1.030 ;
        RECT  7.215 0.630 7.555 1.410 ;
        RECT  7.130 1.180 8.760 1.410 ;
        RECT  9.505 0.800 9.735 1.845 ;
        RECT  9.505 1.615 11.105 1.845 ;
        RECT  10.765 1.615 11.105 1.950 ;
        RECT  8.530 0.800 8.760 2.120 ;
        RECT  8.420 1.780 8.760 2.120 ;
        RECT  7.130 1.180 7.415 2.165 ;
        RECT  7.065 1.825 7.415 2.165 ;
        RECT  7.185 1.180 7.415 2.825 ;
        RECT  7.185 2.540 7.610 2.825 ;
        RECT  8.990 1.260 9.275 1.600 ;
        RECT  6.040 1.760 6.380 2.110 ;
        RECT  6.040 1.880 6.780 2.110 ;
        RECT  10.040 2.175 10.380 2.515 ;
        RECT  10.040 2.280 11.425 2.515 ;
        RECT  9.045 2.285 11.425 2.515 ;
        RECT  11.140 2.280 11.425 2.620 ;
        RECT  6.550 1.880 6.780 3.285 ;
        RECT  8.790 2.805 9.275 3.145 ;
        RECT  9.045 1.260 9.275 3.145 ;
        RECT  6.550 3.055 9.035 3.285 ;
        RECT  11.035 1.090 11.810 1.385 ;
        RECT  11.580 1.090 11.810 2.055 ;
        RECT  11.655 1.835 11.885 3.090 ;
        RECT  13.415 2.750 13.755 3.090 ;
        RECT  10.480 2.860 13.755 3.090 ;
        RECT  10.480 2.860 10.820 3.615 ;
        RECT  12.040 1.320 12.325 1.660 ;
        RECT  12.040 1.430 13.875 1.660 ;
        RECT  13.535 1.430 13.875 2.110 ;
        RECT  13.535 1.880 14.395 2.110 ;
        RECT  13.985 1.880 14.395 2.220 ;
        RECT  13.985 1.880 14.215 3.610 ;
        RECT  13.130 3.380 14.215 3.610 ;
        RECT  13.130 3.380 13.470 3.720 ;
        RECT  1.770 0.940 4.60 1.170 ;
        RECT  2.120 3.500 3.30 3.730 ;
        RECT  9.045 2.285 10.20 2.515 ;
        RECT  6.550 3.055 8.40 3.285 ;
        RECT  10.480 2.860 12.80 3.090 ;
    END
END SDFFSX2

MACRO SDFFSX1
    CLASS CORE ;
    FOREIGN SDFFSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.850 2.860 16.255 3.240 ;
        RECT  15.850 0.940 16.190 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.165 1.640 15.620 2.020 ;
        RECT  14.520 2.870 15.395 3.100 ;
        RECT  15.165 1.235 15.395 3.100 ;
        RECT  14.570 1.235 15.395 1.465 ;
        RECT  14.570 0.700 14.800 1.465 ;
        RECT  14.410 3.625 14.750 3.965 ;
        RECT  14.520 2.870 14.750 3.965 ;
        RECT  14.410 0.700 14.800 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.670 3.995 2.030 4.250 ;
        RECT  1.670 3.960 2.015 4.250 ;
        RECT  1.670 3.470 1.900 4.250 ;
        RECT  1.410 3.470 1.900 3.815 ;
        RECT  1.385 3.470 1.900 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.940 2.800 3.655 3.190 ;
        RECT  2.940 2.045 3.170 3.190 ;
        RECT  0.575 2.045 3.170 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.805 2.710 3.190 ;
        RECT  2.370 2.505 2.710 3.190 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.075 2.250 13.735 2.700 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.265 1.660 8.755 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.130 -0.400 15.470 1.005 ;
        RECT  12.755 -0.400 13.095 1.025 ;
        RECT  10.770 -0.400 11.110 1.005 ;
        RECT  8.705 -0.400 9.045 0.970 ;
        RECT  5.170 -0.400 5.510 0.710 ;
        RECT  2.825 1.090 3.825 1.325 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.130 3.330 15.470 5.280 ;
        RECT  13.825 4.170 14.165 5.280 ;
        RECT  12.330 3.630 12.645 5.280 ;
        RECT  9.765 3.480 10.105 5.280 ;
        RECT  8.465 3.535 8.805 5.280 ;
        RECT  5.170 3.430 5.510 5.280 ;
        RECT  3.470 4.170 3.810 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.690 1.815 ;
        RECT  3.350 1.555 3.690 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  4.080 1.570 4.420 2.090 ;
        RECT  3.920 1.860 5.830 2.090 ;
        RECT  5.490 1.860 5.830 2.280 ;
        RECT  3.920 1.860 4.150 3.190 ;
        RECT  3.920 2.850 4.480 3.190 ;
        RECT  6.325 1.200 6.740 1.540 ;
        RECT  4.390 2.320 4.995 2.605 ;
        RECT  4.780 2.510 6.555 2.740 ;
        RECT  6.325 1.200 6.555 3.385 ;
        RECT  6.325 3.045 6.745 3.385 ;
        RECT  4.710 2.970 5.975 3.200 ;
        RECT  5.745 2.970 5.975 3.845 ;
        RECT  4.710 2.970 4.940 3.650 ;
        RECT  2.130 3.420 4.940 3.650 ;
        RECT  2.130 3.420 2.470 3.760 ;
        RECT  7.165 3.535 7.505 3.845 ;
        RECT  5.745 3.615 7.505 3.845 ;
        RECT  2.255 0.630 4.625 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  4.395 0.630 4.625 1.170 ;
        RECT  5.750 0.740 7.465 0.970 ;
        RECT  4.395 0.940 5.980 1.170 ;
        RECT  7.235 0.740 7.465 1.600 ;
        RECT  7.235 1.260 7.575 1.600 ;
        RECT  9.735 1.240 10.075 1.580 ;
        RECT  9.735 1.240 9.965 3.120 ;
        RECT  6.785 1.770 7.070 2.700 ;
        RECT  8.350 2.625 9.965 2.965 ;
        RECT  6.975 2.470 7.205 3.305 ;
        RECT  9.735 2.890 11.020 3.120 ;
        RECT  10.680 2.890 11.020 3.230 ;
        RECT  8.350 2.625 8.580 3.305 ;
        RECT  6.975 3.075 8.580 3.305 ;
        RECT  9.275 0.780 10.540 1.010 ;
        RECT  7.805 0.630 8.245 1.430 ;
        RECT  9.275 0.780 9.505 1.430 ;
        RECT  7.805 1.200 9.505 1.430 ;
        RECT  8.985 1.200 9.215 2.105 ;
        RECT  8.985 1.765 9.325 2.105 ;
        RECT  7.805 0.630 8.035 2.235 ;
        RECT  7.400 1.950 8.005 2.290 ;
        RECT  10.310 2.220 10.825 2.450 ;
        RECT  10.310 0.780 10.540 2.450 ;
        RECT  10.485 2.330 11.640 2.560 ;
        RECT  7.665 1.950 8.005 2.845 ;
        RECT  11.355 2.330 11.640 3.450 ;
        RECT  13.510 0.670 13.850 1.010 ;
        RECT  13.510 0.670 13.740 1.485 ;
        RECT  11.525 1.255 13.740 1.485 ;
        RECT  11.525 1.255 12.100 1.610 ;
        RECT  11.870 1.255 12.100 3.970 ;
        RECT  10.960 3.680 12.100 3.970 ;
        RECT  14.030 1.640 14.370 2.640 ;
        RECT  14.030 2.300 14.780 2.640 ;
        RECT  12.330 2.645 12.670 3.160 ;
        RECT  14.030 1.640 14.260 3.160 ;
        RECT  12.330 2.930 14.260 3.160 ;
        RECT  13.025 2.930 13.365 3.970 ;
        RECT  1.255 1.585 2.40 1.815 ;
        RECT  2.130 3.420 3.90 3.650 ;
        RECT  2.255 0.630 3.50 0.860 ;
        RECT  11.525 1.255 12.60 1.485 ;
    END
END SDFFSX1

MACRO SDFFSX0
    CLASS CORE ;
    FOREIGN SDFFSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.480 2.640 14.995 3.240 ;
        RECT  14.670 1.170 14.995 3.240 ;
        RECT  14.560 1.170 14.995 1.510 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.610  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 1.640 14.365 2.020 ;
        RECT  13.590 2.620 14.215 2.960 ;
        RECT  13.985 0.630 14.215 2.960 ;
        RECT  13.305 0.630 14.215 0.890 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 2.250 12.690 2.660 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.675 2.230 8.175 2.695 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.480 3.470 14.820 5.280 ;
        RECT  13.190 4.165 13.530 5.280 ;
        RECT  11.715 3.630 12.000 5.280 ;
        RECT  8.960 3.630 9.300 5.280 ;
        RECT  8.025 3.880 8.365 5.280 ;
        RECT  4.830 3.910 5.115 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  14.560 -0.400 14.900 0.710 ;
        RECT  12.195 -0.400 12.535 0.890 ;
        RECT  10.110 -0.400 10.395 0.710 ;
        RECT  10.090 -0.400 10.395 0.675 ;
        RECT  8.165 -0.400 8.500 1.030 ;
        RECT  4.495 -0.400 4.835 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.815 ;
        RECT  2.930 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.505 1.805 5.295 2.035 ;
        RECT  3.505 1.805 3.970 2.095 ;
        RECT  5.010 1.805 5.295 2.205 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.525 1.230 6.430 1.540 ;
        RECT  3.965 2.325 4.250 2.665 ;
        RECT  3.965 2.435 5.755 2.665 ;
        RECT  5.525 1.230 5.755 3.220 ;
        RECT  5.520 2.435 5.755 3.220 ;
        RECT  5.520 2.990 6.235 3.220 ;
        RECT  6.005 2.990 6.235 3.790 ;
        RECT  6.005 3.450 6.345 3.790 ;
        RECT  4.370 3.450 5.575 3.680 ;
        RECT  4.370 3.450 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.345 3.450 5.575 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.765 3.880 7.105 4.250 ;
        RECT  5.345 4.020 7.105 4.250 ;
        RECT  5.065 0.770 7.255 1.000 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  5.065 0.770 5.295 1.355 ;
        RECT  1.980 1.125 5.295 1.355 ;
        RECT  6.915 0.770 7.255 1.540 ;
        RECT  5.985 2.440 6.325 2.760 ;
        RECT  5.985 2.530 6.805 2.760 ;
        RECT  9.190 1.230 9.420 3.245 ;
        RECT  8.625 2.905 10.250 3.245 ;
        RECT  9.190 2.850 10.250 3.245 ;
        RECT  7.795 3.015 10.250 3.245 ;
        RECT  6.575 2.530 6.805 3.650 ;
        RECT  7.795 3.015 8.025 3.650 ;
        RECT  6.575 3.420 8.025 3.650 ;
        RECT  8.730 0.770 9.880 1.000 ;
        RECT  8.730 0.770 8.960 1.590 ;
        RECT  7.615 1.360 8.960 1.590 ;
        RECT  7.615 1.360 7.955 2.000 ;
        RECT  5.985 1.770 7.955 2.000 ;
        RECT  9.650 0.770 9.880 2.290 ;
        RECT  5.985 1.770 7.445 2.110 ;
        RECT  8.565 1.360 8.905 2.160 ;
        RECT  9.650 2.060 10.265 2.290 ;
        RECT  9.925 2.170 10.935 2.400 ;
        RECT  7.215 1.770 7.445 3.190 ;
        RECT  7.215 2.880 7.530 3.190 ;
        RECT  10.705 2.170 10.935 3.440 ;
        RECT  7.215 2.905 7.565 3.190 ;
        RECT  10.705 3.100 10.975 3.440 ;
        RECT  10.965 1.110 11.505 1.450 ;
        RECT  11.210 1.110 11.505 3.385 ;
        RECT  12.540 3.045 12.860 3.385 ;
        RECT  11.210 3.155 12.860 3.385 ;
        RECT  11.210 1.110 11.440 3.970 ;
        RECT  10.255 3.670 11.440 3.970 ;
        RECT  13.305 1.315 13.645 2.320 ;
        RECT  11.925 1.700 13.645 2.020 ;
        RECT  13.090 1.980 13.755 2.320 ;
        RECT  13.090 1.700 13.320 3.900 ;
        RECT  12.390 3.650 13.320 3.900 ;
        RECT  12.390 3.650 12.730 3.970 ;
        RECT  0.980 1.585 2.80 1.815 ;
        RECT  1.995 3.710 3.50 3.940 ;
        RECT  5.065 0.770 6.70 1.000 ;
        RECT  1.980 1.125 4.70 1.355 ;
        RECT  7.795 3.015 9.30 3.245 ;
    END
END SDFFSX0

MACRO SDFFSQX4
    CLASS CORE ;
    FOREIGN SDFFSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.075 2.250 17.415 4.100 ;
        RECT  15.635 2.250 17.415 2.630 ;
        RECT  16.560 1.230 16.900 2.630 ;
        RECT  15.635 2.250 15.975 4.100 ;
        RECT  15.540 0.700 15.770 2.480 ;
        RECT  15.240 0.700 15.770 1.040 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.760 1.640 14.365 2.020 ;
        RECT  13.760 1.640 14.105 2.200 ;
        END
    END SN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 1.640 8.920 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  17.120 -0.400 17.460 0.710 ;
        RECT  16.000 -0.400 16.340 0.710 ;
        RECT  13.190 -0.400 14.000 0.800 ;
        RECT  10.715 -0.400 11.000 1.370 ;
        RECT  8.820 -0.400 9.105 0.950 ;
        RECT  3.400 -0.400 5.150 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.355 2.860 16.695 5.280 ;
        RECT  14.875 4.140 15.215 5.280 ;
        RECT  13.590 2.890 13.930 5.280 ;
        RECT  11.370 3.965 11.710 5.280 ;
        RECT  8.975 2.910 9.260 5.280 ;
        RECT  4.795 3.965 5.135 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.585 5.740 1.875 ;
        RECT  5.400 1.585 5.740 2.265 ;
        RECT  3.895 1.585 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.025 1.190 6.800 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  6.025 1.190 6.255 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  6.025 2.935 6.450 3.275 ;
        RECT  4.630 3.045 6.450 3.275 ;
        RECT  6.830 2.980 7.165 3.735 ;
        RECT  2.020 3.505 7.165 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.380 0.730 7.260 0.960 ;
        RECT  2.255 0.940 5.610 1.170 ;
        RECT  7.030 0.730 7.260 1.660 ;
        RECT  7.030 1.320 7.615 1.660 ;
        RECT  9.335 0.775 10.485 1.005 ;
        RECT  7.490 0.735 8.360 1.090 ;
        RECT  7.855 0.735 8.360 1.410 ;
        RECT  7.855 1.180 9.565 1.410 ;
        RECT  10.255 0.775 10.485 1.960 ;
        RECT  10.255 1.730 11.910 1.960 ;
        RECT  11.570 1.730 11.910 2.070 ;
        RECT  9.335 0.775 9.565 2.100 ;
        RECT  9.210 1.760 9.565 2.100 ;
        RECT  7.855 0.735 8.085 2.940 ;
        RECT  7.855 2.600 8.285 2.940 ;
        RECT  6.485 1.840 6.795 2.195 ;
        RECT  6.485 1.965 7.625 2.195 ;
        RECT  9.795 1.240 10.025 2.680 ;
        RECT  9.795 2.340 10.740 2.680 ;
        RECT  12.240 1.540 12.525 2.680 ;
        RECT  8.515 2.450 12.525 2.680 ;
        RECT  9.640 2.450 9.980 2.860 ;
        RECT  7.395 1.965 7.625 3.400 ;
        RECT  8.515 2.450 8.745 3.400 ;
        RECT  7.395 3.170 8.745 3.400 ;
        RECT  9.640 2.450 9.870 3.855 ;
        RECT  10.840 3.505 12.180 3.735 ;
        RECT  11.950 3.505 12.180 4.100 ;
        RECT  9.640 3.625 11.070 3.855 ;
        RECT  11.950 3.760 12.460 4.100 ;
        RECT  11.810 0.970 12.150 1.310 ;
        RECT  11.810 1.080 12.985 1.310 ;
        RECT  14.505 2.320 14.845 2.660 ;
        RECT  12.755 2.430 14.845 2.660 ;
        RECT  12.755 1.080 12.985 3.220 ;
        RECT  10.180 2.990 12.985 3.220 ;
        RECT  12.360 2.990 12.700 3.330 ;
        RECT  10.180 2.990 10.520 3.395 ;
        RECT  13.215 1.180 15.010 1.410 ;
        RECT  14.670 1.180 15.010 1.700 ;
        RECT  13.215 1.180 13.500 1.530 ;
        RECT  14.670 1.470 15.310 1.700 ;
        RECT  15.080 1.470 15.310 3.120 ;
        RECT  14.315 2.890 15.310 3.120 ;
        RECT  14.315 2.890 14.655 3.730 ;
        RECT  1.145 1.585 2.20 1.815 ;
        RECT  2.020 3.505 6.60 3.735 ;
        RECT  2.255 0.940 4.80 1.170 ;
        RECT  8.515 2.450 11.90 2.680 ;
        RECT  12.755 2.430 13.50 2.660 ;
        RECT  10.180 2.990 11.60 3.220 ;
    END
END SDFFSQX4

MACRO SDFFSQX2
    CLASS CORE ;
    FOREIGN SDFFSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.670 1.250 15.010 2.630 ;
        RECT  14.450 2.250 14.790 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.720 1.005 2.200 ;
        END
    END SE
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.585 2.050 13.105 2.630 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.645 1.640 8.115 2.160 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.230 -0.400 15.570 0.720 ;
        RECT  14.110 -0.400 14.450 0.720 ;
        RECT  12.300 -0.400 12.645 1.090 ;
        RECT  9.975 -0.400 10.315 0.710 ;
        RECT  8.015 -0.400 8.300 0.950 ;
        RECT  4.530 -0.400 4.870 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.210 3.270 15.550 5.280 ;
        RECT  13.690 4.170 14.030 5.280 ;
        RECT  12.410 3.385 12.750 5.280 ;
        RECT  11.710 3.375 12.050 5.280 ;
        RECT  9.330 3.480 9.670 5.280 ;
        RECT  8.030 3.515 8.370 5.280 ;
        RECT  4.715 3.900 5.055 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.330 2.015 ;
        RECT  4.990 1.785 5.330 2.470 ;
        RECT  3.480 1.400 3.710 3.270 ;
        RECT  3.480 2.930 4.250 3.265 ;
        RECT  3.480 2.930 4.240 3.270 ;
        RECT  5.580 1.190 6.100 1.530 ;
        RECT  3.940 2.245 4.715 2.585 ;
        RECT  4.485 2.245 4.715 2.930 ;
        RECT  5.580 1.190 5.810 3.210 ;
        RECT  4.485 2.700 5.810 2.930 ;
        RECT  5.580 2.870 6.285 3.210 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  5.120 0.730 6.900 0.960 ;
        RECT  1.770 0.940 5.350 1.170 ;
        RECT  6.560 0.730 6.900 1.595 ;
        RECT  4.400 3.440 5.525 3.670 ;
        RECT  2.120 3.500 4.560 3.730 ;
        RECT  5.295 3.515 7.045 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  8.530 0.800 9.735 1.030 ;
        RECT  7.215 0.630 7.555 1.410 ;
        RECT  7.130 1.180 8.760 1.410 ;
        RECT  9.505 0.800 9.735 1.845 ;
        RECT  9.505 1.615 11.105 1.845 ;
        RECT  10.765 1.615 11.105 1.950 ;
        RECT  8.530 0.800 8.760 2.120 ;
        RECT  8.420 1.780 8.760 2.120 ;
        RECT  7.130 1.180 7.415 2.165 ;
        RECT  7.065 1.825 7.415 2.165 ;
        RECT  7.185 1.180 7.415 2.825 ;
        RECT  7.185 2.540 7.610 2.825 ;
        RECT  8.990 1.260 9.275 1.600 ;
        RECT  6.040 1.760 6.380 2.110 ;
        RECT  6.040 1.880 6.780 2.110 ;
        RECT  10.040 2.175 10.380 2.515 ;
        RECT  10.040 2.280 11.425 2.515 ;
        RECT  9.045 2.285 11.425 2.515 ;
        RECT  11.140 2.280 11.425 2.620 ;
        RECT  6.550 1.880 6.780 3.285 ;
        RECT  8.790 2.805 9.275 3.145 ;
        RECT  9.045 1.260 9.275 3.145 ;
        RECT  6.550 3.055 9.035 3.285 ;
        RECT  11.035 1.090 11.810 1.385 ;
        RECT  11.580 1.090 11.810 2.055 ;
        RECT  11.655 1.835 11.885 3.090 ;
        RECT  13.415 2.750 13.755 3.090 ;
        RECT  10.480 2.860 13.755 3.090 ;
        RECT  10.480 2.860 10.820 3.615 ;
        RECT  13.335 0.630 13.675 1.660 ;
        RECT  12.040 1.320 13.675 1.660 ;
        RECT  12.040 1.430 14.215 1.660 ;
        RECT  13.985 1.430 14.215 3.720 ;
        RECT  13.130 3.380 14.215 3.720 ;
        RECT  1.770 0.940 4.70 1.170 ;
        RECT  2.120 3.500 3.60 3.730 ;
        RECT  9.045 2.285 10.90 2.515 ;
        RECT  6.550 3.055 8.70 3.285 ;
        RECT  10.480 2.860 12.60 3.090 ;
        RECT  12.040 1.430 13.70 1.660 ;
    END
END SDFFSQX2

MACRO SDFFSQX1
    CLASS CORE ;
    FOREIGN SDFFSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.250 14.995 2.630 ;
        RECT  14.410 3.625 14.845 3.965 ;
        RECT  14.615 0.700 14.845 3.965 ;
        RECT  14.410 0.700 14.845 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.670 3.995 2.030 4.250 ;
        RECT  1.670 3.960 2.015 4.250 ;
        RECT  1.670 3.470 1.900 4.250 ;
        RECT  1.410 3.470 1.900 3.815 ;
        RECT  1.385 3.470 1.900 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.940 2.800 3.655 3.190 ;
        RECT  2.940 2.045 3.170 3.190 ;
        RECT  0.575 2.045 3.170 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.805 2.710 3.190 ;
        RECT  2.370 2.505 2.710 3.190 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.075 2.250 13.735 2.700 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.265 1.660 8.755 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.130 -0.400 15.470 1.060 ;
        RECT  12.755 -0.400 13.095 1.025 ;
        RECT  10.770 -0.400 11.110 1.005 ;
        RECT  8.705 -0.400 9.045 0.970 ;
        RECT  5.170 -0.400 5.510 0.710 ;
        RECT  2.825 1.090 3.825 1.325 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.130 3.330 15.470 5.280 ;
        RECT  13.825 4.170 14.165 5.280 ;
        RECT  12.330 3.630 12.645 5.280 ;
        RECT  9.765 3.480 10.105 5.280 ;
        RECT  8.465 3.535 8.805 5.280 ;
        RECT  5.170 3.430 5.510 5.280 ;
        RECT  3.470 4.170 3.810 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.690 1.815 ;
        RECT  3.350 1.555 3.690 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  4.080 1.570 4.420 2.090 ;
        RECT  3.920 1.860 5.830 2.090 ;
        RECT  5.490 1.860 5.830 2.280 ;
        RECT  3.920 1.860 4.150 3.190 ;
        RECT  3.920 2.850 4.480 3.190 ;
        RECT  6.325 1.200 6.740 1.540 ;
        RECT  4.390 2.320 4.995 2.605 ;
        RECT  4.780 2.510 6.555 2.740 ;
        RECT  6.325 1.200 6.555 3.385 ;
        RECT  6.325 3.045 6.745 3.385 ;
        RECT  4.710 2.970 5.975 3.200 ;
        RECT  5.745 2.970 5.975 3.845 ;
        RECT  4.710 2.970 4.940 3.650 ;
        RECT  2.130 3.420 4.940 3.650 ;
        RECT  2.130 3.420 2.470 3.760 ;
        RECT  7.165 3.535 7.505 3.845 ;
        RECT  5.745 3.615 7.505 3.845 ;
        RECT  2.255 0.630 4.625 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  4.395 0.630 4.625 1.170 ;
        RECT  5.750 0.740 7.465 0.970 ;
        RECT  4.395 0.940 5.980 1.170 ;
        RECT  7.235 0.740 7.465 1.600 ;
        RECT  7.235 1.260 7.575 1.600 ;
        RECT  9.735 1.240 10.075 1.580 ;
        RECT  9.735 1.240 9.965 3.120 ;
        RECT  6.785 1.770 7.070 2.700 ;
        RECT  8.350 2.625 9.965 2.965 ;
        RECT  6.975 2.470 7.205 3.305 ;
        RECT  9.735 2.890 11.020 3.120 ;
        RECT  10.680 2.890 11.020 3.230 ;
        RECT  8.350 2.625 8.580 3.305 ;
        RECT  6.975 3.075 8.580 3.305 ;
        RECT  9.275 0.780 10.540 1.010 ;
        RECT  7.805 0.630 8.245 1.430 ;
        RECT  9.275 0.780 9.505 1.430 ;
        RECT  7.805 1.200 9.505 1.430 ;
        RECT  8.985 1.200 9.215 2.105 ;
        RECT  8.985 1.765 9.325 2.105 ;
        RECT  7.805 0.630 8.035 2.235 ;
        RECT  7.400 1.950 8.005 2.290 ;
        RECT  10.310 2.220 10.825 2.450 ;
        RECT  10.310 0.780 10.540 2.450 ;
        RECT  10.485 2.330 11.640 2.560 ;
        RECT  7.665 1.950 8.005 2.845 ;
        RECT  11.355 2.330 11.640 3.450 ;
        RECT  13.510 0.910 13.850 1.250 ;
        RECT  13.510 0.910 13.740 1.485 ;
        RECT  11.525 1.255 13.740 1.485 ;
        RECT  11.525 1.255 12.100 1.610 ;
        RECT  11.870 1.255 12.100 3.970 ;
        RECT  10.960 3.680 12.100 3.970 ;
        RECT  14.030 1.640 14.370 1.980 ;
        RECT  12.330 2.645 12.670 3.160 ;
        RECT  14.030 1.640 14.260 3.160 ;
        RECT  12.330 2.930 14.260 3.160 ;
        RECT  13.025 2.930 13.365 3.970 ;
        RECT  1.255 1.585 2.60 1.815 ;
        RECT  2.130 3.420 3.80 3.650 ;
        RECT  2.255 0.630 3.30 0.860 ;
        RECT  11.525 1.255 12.40 1.485 ;
    END
END SDFFSQX1

MACRO SDFFSQX0
    CLASS CORE ;
    FOREIGN SDFFSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.595  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.340 2.250 13.745 2.980 ;
        RECT  13.515 0.630 13.745 2.980 ;
        RECT  12.990 0.630 13.745 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.980 2.240 12.585 2.705 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 2.170 8.115 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.940 4.165 13.280 5.280 ;
        RECT  11.395 3.910 11.680 5.280 ;
        RECT  8.760 3.630 9.100 5.280 ;
        RECT  8.025 3.880 8.365 5.280 ;
        RECT  4.830 3.910 5.115 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  11.880 -0.400 12.220 0.910 ;
        RECT  9.850 -0.400 10.190 0.710 ;
        RECT  7.900 -0.400 8.185 0.970 ;
        RECT  4.495 -0.400 4.835 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.505 1.805 5.295 2.095 ;
        RECT  5.010 1.805 5.295 2.205 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.525 1.230 6.430 1.540 ;
        RECT  3.965 2.325 4.250 2.665 ;
        RECT  3.965 2.435 5.755 2.665 ;
        RECT  5.525 1.230 5.755 3.220 ;
        RECT  5.520 2.435 5.755 3.220 ;
        RECT  5.520 2.990 6.235 3.220 ;
        RECT  6.005 2.990 6.235 3.790 ;
        RECT  6.005 3.450 6.345 3.790 ;
        RECT  4.370 3.450 5.575 3.680 ;
        RECT  4.370 3.450 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.345 3.450 5.575 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.765 3.880 7.105 4.250 ;
        RECT  5.345 4.020 7.105 4.250 ;
        RECT  5.065 0.630 7.110 0.860 ;
        RECT  6.770 0.630 7.110 0.970 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  5.065 0.630 5.295 1.355 ;
        RECT  1.980 1.125 5.295 1.355 ;
        RECT  8.875 1.230 9.160 1.570 ;
        RECT  5.985 2.440 6.325 2.760 ;
        RECT  5.985 2.530 6.805 2.760 ;
        RECT  8.930 2.710 10.050 2.940 ;
        RECT  9.710 2.600 10.050 2.940 ;
        RECT  8.930 1.230 9.160 3.220 ;
        RECT  8.300 2.890 9.160 3.220 ;
        RECT  6.575 2.530 6.805 3.650 ;
        RECT  8.300 2.890 8.530 3.650 ;
        RECT  6.575 3.420 8.530 3.650 ;
        RECT  8.415 0.770 9.620 1.000 ;
        RECT  7.105 1.250 8.645 1.490 ;
        RECT  7.105 1.250 7.730 1.535 ;
        RECT  8.415 0.770 8.645 2.110 ;
        RECT  8.345 1.250 8.645 2.110 ;
        RECT  9.390 0.770 9.620 2.160 ;
        RECT  7.105 1.250 7.440 2.110 ;
        RECT  5.985 1.770 7.440 2.110 ;
        RECT  8.345 1.770 8.685 2.110 ;
        RECT  9.390 1.930 10.265 2.160 ;
        RECT  9.925 2.040 10.595 2.270 ;
        RECT  7.210 1.250 7.440 3.190 ;
        RECT  10.365 2.040 10.595 3.415 ;
        RECT  7.210 2.850 7.565 3.190 ;
        RECT  10.365 3.075 10.705 3.415 ;
        RECT  10.650 1.110 11.165 1.450 ;
        RECT  10.935 2.990 12.630 3.330 ;
        RECT  10.935 1.110 11.165 3.970 ;
        RECT  9.990 3.645 11.165 3.970 ;
        RECT  12.990 1.350 13.285 1.915 ;
        RECT  11.610 1.700 13.090 2.010 ;
        RECT  12.860 1.700 13.090 3.790 ;
        RECT  12.140 3.560 13.090 3.790 ;
        RECT  12.140 3.560 12.480 3.880 ;
        RECT  0.980 1.585 2.60 1.960 ;
        RECT  1.995 3.710 3.70 3.940 ;
        RECT  5.065 0.630 6.60 0.860 ;
        RECT  1.980 1.125 4.60 1.355 ;
    END
END SDFFSQX0

MACRO SDFFRX4
    CLASS CORE ;
    FOREIGN SDFFRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.050 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  21.530 1.130 21.870 4.005 ;
        RECT  20.090 2.250 21.870 2.630 ;
        RECT  20.090 1.130 20.430 4.005 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.119  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.355 3.010 19.730 3.240 ;
        RECT  19.500 1.700 19.730 3.240 ;
        RECT  17.210 1.700 19.730 1.930 ;
        RECT  18.795 3.010 19.135 3.350 ;
        RECT  18.650 1.130 18.990 1.930 ;
        RECT  17.355 2.860 18.145 3.240 ;
        RECT  17.355 2.860 17.695 4.130 ;
        RECT  17.210 1.130 17.550 1.930 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.020 1.640 15.650 2.175 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.660 10.630 2.135 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 22.050 0.400 ;
        RECT  20.810 -0.400 21.150 1.470 ;
        RECT  19.370 -0.400 19.710 1.470 ;
        RECT  17.930 -0.400 18.270 1.470 ;
        RECT  15.670 -0.400 16.010 0.950 ;
        RECT  9.920 -0.400 10.205 0.970 ;
        RECT  4.775 -0.400 5.915 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 22.050 5.280 ;
        RECT  20.810 2.860 21.150 5.280 ;
        RECT  19.370 3.665 19.710 5.280 ;
        RECT  18.075 3.470 18.415 5.280 ;
        RECT  16.595 4.170 16.935 5.280 ;
        RECT  14.155 3.640 15.615 5.280 ;
        RECT  11.745 3.980 12.085 5.280 ;
        RECT  9.135 2.950 9.475 5.280 ;
        RECT  4.660 4.115 5.700 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 5.885 2.095 ;
        RECT  5.655 1.860 5.885 2.800 ;
        RECT  5.655 2.460 5.995 2.800 ;
        RECT  3.895 1.815 4.125 3.425 ;
        RECT  3.895 3.085 4.260 3.425 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 6.625 1.585 ;
        RECT  5.015 1.355 6.625 1.630 ;
        RECT  6.335 1.355 6.625 1.695 ;
        RECT  7.530 3.020 7.870 3.360 ;
        RECT  2.020 3.655 6.390 3.885 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  7.530 3.020 7.760 4.000 ;
        RECT  6.160 3.770 7.760 4.000 ;
        RECT  6.855 1.160 7.900 1.500 ;
        RECT  4.355 2.325 4.640 2.665 ;
        RECT  4.355 2.435 4.890 2.665 ;
        RECT  4.660 2.435 4.890 3.425 ;
        RECT  4.660 3.085 5.000 3.425 ;
        RECT  4.660 3.195 7.085 3.425 ;
        RECT  6.855 1.160 7.085 3.450 ;
        RECT  6.745 3.110 7.085 3.450 ;
        RECT  6.210 0.630 8.360 0.860 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.210 0.630 6.440 1.125 ;
        RECT  4.315 0.895 6.440 1.125 ;
        RECT  8.130 0.630 8.360 1.660 ;
        RECT  8.130 1.320 8.715 1.660 ;
        RECT  8.920 2.395 9.260 2.680 ;
        RECT  10.895 1.240 11.125 2.680 ;
        RECT  8.920 2.450 11.125 2.680 ;
        RECT  9.855 2.450 10.195 3.915 ;
        RECT  11.215 3.520 12.545 3.750 ;
        RECT  12.315 3.520 12.545 4.130 ;
        RECT  9.855 3.685 11.445 3.915 ;
        RECT  12.315 3.790 13.545 4.130 ;
        RECT  10.435 0.775 11.585 1.005 ;
        RECT  9.120 0.735 9.460 1.090 ;
        RECT  10.435 0.775 10.665 1.430 ;
        RECT  9.230 1.200 10.665 1.430 ;
        RECT  7.315 1.810 7.655 2.150 ;
        RECT  11.355 0.775 11.585 2.185 ;
        RECT  9.230 0.735 9.460 2.150 ;
        RECT  7.315 1.920 9.460 2.150 ;
        RECT  13.350 1.555 13.690 2.185 ;
        RECT  11.355 1.955 13.690 2.185 ;
        RECT  12.495 1.955 12.835 2.755 ;
        RECT  8.350 1.920 8.690 3.860 ;
        RECT  11.815 0.630 15.210 0.860 ;
        RECT  14.385 0.630 15.210 0.950 ;
        RECT  11.815 0.630 12.110 1.500 ;
        RECT  12.920 1.090 14.150 1.320 ;
        RECT  15.950 2.370 16.290 2.710 ;
        RECT  13.920 2.480 16.290 2.710 ;
        RECT  14.715 2.480 15.055 3.050 ;
        RECT  13.920 1.090 14.150 3.215 ;
        RECT  10.555 2.985 14.150 3.215 ;
        RECT  12.795 2.985 13.135 3.450 ;
        RECT  10.555 2.985 10.895 3.455 ;
        RECT  14.380 1.180 16.770 1.410 ;
        RECT  16.430 1.180 16.770 1.520 ;
        RECT  14.380 1.180 14.720 1.680 ;
        RECT  16.540 2.310 19.270 2.540 ;
        RECT  18.985 2.310 19.270 2.650 ;
        RECT  16.540 1.180 16.770 3.170 ;
        RECT  16.035 2.940 16.770 3.170 ;
        RECT  16.035 2.940 16.375 3.760 ;
        RECT  1.145 1.585 2.90 1.815 ;
        RECT  1.605 1.125 3.70 1.355 ;
        RECT  3.855 1.355 5.00 1.585 ;
        RECT  2.020 3.655 5.30 3.885 ;
        RECT  4.660 3.195 6.20 3.425 ;
        RECT  6.210 0.630 7.70 0.860 ;
        RECT  2.255 0.630 3.70 0.895 ;
        RECT  4.315 0.895 5.60 1.125 ;
        RECT  8.920 2.450 10.50 2.680 ;
        RECT  7.315 1.920 8.80 2.150 ;
        RECT  11.355 1.955 12.20 2.185 ;
        RECT  11.815 0.630 14.30 0.860 ;
        RECT  13.920 2.480 15.20 2.710 ;
        RECT  10.555 2.985 13.50 3.215 ;
        RECT  14.380 1.180 15.10 1.410 ;
        RECT  16.540 2.310 18.40 2.540 ;
    END
END SDFFRX4

MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.270 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.020 0.820 16.255 3.240 ;
        RECT  15.710 2.860 16.105 3.830 ;
        RECT  15.870 0.820 16.255 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.200 2.110 13.735 2.675 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.135 1.230 17.530 2.020 ;
        RECT  17.030 2.640 17.370 3.550 ;
        RECT  17.135 1.230 17.370 3.550 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.250 9.630 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.270 0.400 ;
        RECT  17.750 -0.400 18.090 0.710 ;
        RECT  16.630 -0.400 16.970 0.710 ;
        RECT  15.110 -0.400 15.450 0.970 ;
        RECT  14.005 -0.400 14.345 1.220 ;
        RECT  9.035 -0.400 9.320 1.360 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.270 5.280 ;
        RECT  17.750 2.640 18.090 5.280 ;
        RECT  16.470 3.950 16.810 5.280 ;
        RECT  14.950 3.775 15.290 5.280 ;
        RECT  12.745 3.365 13.085 5.280 ;
        RECT  9.895 3.525 10.235 5.280 ;
        RECT  8.595 3.440 8.935 5.280 ;
        RECT  4.655 3.960 5.645 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.685 ;
        RECT  4.710 1.400 5.915 1.685 ;
        RECT  4.135 1.550 4.475 2.180 ;
        RECT  3.895 1.950 6.165 2.180 ;
        RECT  5.825 1.950 6.165 2.375 ;
        RECT  3.895 1.950 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.805 1.260 7.145 1.600 ;
        RECT  6.495 1.370 7.145 1.600 ;
        RECT  4.415 2.410 5.045 2.750 ;
        RECT  4.705 2.410 5.045 3.270 ;
        RECT  6.495 1.370 6.725 3.270 ;
        RECT  4.705 3.040 6.875 3.270 ;
        RECT  6.535 3.040 6.875 3.625 ;
        RECT  2.120 3.500 6.305 3.730 ;
        RECT  6.075 3.500 6.305 4.125 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  7.295 3.535 7.635 4.125 ;
        RECT  6.075 3.895 7.635 4.125 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.800 7.945 1.030 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  7.605 0.800 7.945 1.600 ;
        RECT  8.425 2.305 8.715 3.165 ;
        RECT  10.010 1.260 10.240 3.165 ;
        RECT  8.425 2.860 10.240 3.165 ;
        RECT  8.425 2.935 10.870 3.165 ;
        RECT  10.640 2.935 10.870 4.145 ;
        RECT  10.640 3.915 12.160 4.145 ;
        RECT  11.820 3.915 12.160 4.250 ;
        RECT  9.550 0.800 10.700 1.030 ;
        RECT  9.550 0.800 9.780 1.820 ;
        RECT  8.260 1.590 9.780 1.820 ;
        RECT  8.260 0.630 8.600 2.060 ;
        RECT  6.955 1.830 8.600 2.060 ;
        RECT  6.955 1.830 8.165 2.220 ;
        RECT  10.470 0.800 10.700 2.455 ;
        RECT  10.470 2.225 11.150 2.455 ;
        RECT  11.995 2.225 12.320 2.565 ;
        RECT  10.810 2.330 12.320 2.565 ;
        RECT  7.825 1.830 8.165 3.175 ;
        RECT  10.930 0.630 13.625 0.860 ;
        RECT  13.285 0.630 13.625 1.105 ;
        RECT  10.930 0.630 11.215 1.330 ;
        RECT  12.055 1.090 12.780 1.375 ;
        RECT  13.965 2.400 14.935 2.740 ;
        RECT  12.550 1.090 12.780 3.135 ;
        RECT  13.965 2.400 14.195 3.135 ;
        RECT  11.300 2.905 14.195 3.135 ;
        RECT  11.300 2.905 11.640 3.685 ;
        RECT  13.465 2.905 13.805 4.175 ;
        RECT  13.010 1.380 13.355 1.720 ;
        RECT  13.010 1.490 15.145 1.720 ;
        RECT  14.805 1.490 15.145 2.100 ;
        RECT  14.805 1.870 15.665 2.100 ;
        RECT  15.165 1.870 15.665 2.210 ;
        RECT  15.165 1.870 15.395 3.310 ;
        RECT  14.425 2.970 15.395 3.310 ;
        RECT  1.255 1.585 2.80 1.815 ;
        RECT  2.825 1.090 3.40 1.320 ;
        RECT  1.715 1.125 2.40 1.355 ;
        RECT  3.895 1.950 5.30 2.180 ;
        RECT  4.705 3.040 5.20 3.270 ;
        RECT  2.120 3.500 5.50 3.730 ;
        RECT  2.255 0.630 4.00 0.860 ;
        RECT  8.425 2.935 9.40 3.165 ;
        RECT  10.930 0.630 12.80 0.860 ;
        RECT  11.300 2.905 13.40 3.135 ;
        RECT  13.010 1.490 14.90 1.720 ;
    END
END SDFFRX2

MACRO SDFFRX1
    CLASS CORE ;
    FOREIGN SDFFRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.865 0.940 16.255 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.245 1.640 15.635 2.020 ;
        RECT  14.735 2.870 15.480 3.100 ;
        RECT  15.245 1.640 15.480 3.100 ;
        RECT  15.245 1.260 15.475 3.100 ;
        RECT  14.680 1.260 15.475 1.490 ;
        RECT  14.420 3.780 14.965 4.120 ;
        RECT  14.735 2.870 14.965 4.120 ;
        RECT  14.680 0.700 14.910 1.490 ;
        RECT  14.420 0.700 14.910 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.665 3.995 2.030 4.250 ;
        RECT  1.665 3.960 2.010 4.250 ;
        RECT  1.665 3.470 1.895 4.250 ;
        RECT  1.410 3.470 1.895 3.815 ;
        RECT  1.385 3.470 1.895 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.970 2.800 3.655 3.240 ;
        RECT  2.970 2.045 3.200 3.240 ;
        RECT  0.575 2.045 3.200 2.275 ;
        RECT  0.575 1.660 0.860 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.745 2.170 13.280 2.630 ;
        END
    END RN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.030 1.660 9.480 2.130 ;
        RECT  8.945 1.660 9.480 2.030 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.140 -0.400 15.480 1.030 ;
        RECT  13.460 -0.400 13.800 0.975 ;
        RECT  8.820 -0.400 9.105 0.970 ;
        RECT  4.815 -0.400 5.155 0.655 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.195 3.330 15.480 5.280 ;
        RECT  12.740 3.820 13.085 5.280 ;
        RECT  10.125 3.470 10.465 5.280 ;
        RECT  8.825 3.160 9.165 5.280 ;
        RECT  4.910 3.845 5.870 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.130 0.900 1.430 ;
        RECT  0.115 1.200 1.485 1.430 ;
        RECT  1.255 1.200 1.485 1.815 ;
        RECT  1.255 1.585 3.665 1.815 ;
        RECT  3.380 1.555 3.665 1.895 ;
        RECT  0.115 1.130 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.125 1.320 ;
        RECT  3.485 1.090 4.125 1.325 ;
        RECT  3.895 1.090 4.125 1.580 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  3.895 1.345 5.685 1.580 ;
        RECT  5.345 1.345 5.685 1.650 ;
        RECT  3.900 1.810 5.170 2.040 ;
        RECT  5.000 1.880 5.965 2.220 ;
        RECT  3.900 1.810 4.220 3.425 ;
        RECT  6.320 1.230 6.915 1.540 ;
        RECT  4.450 2.325 4.760 3.155 ;
        RECT  6.320 1.230 6.550 3.155 ;
        RECT  4.450 2.870 6.550 3.155 ;
        RECT  4.450 2.925 7.100 3.155 ;
        RECT  6.760 2.925 7.100 3.385 ;
        RECT  2.255 0.630 4.585 0.860 ;
        RECT  4.355 0.630 4.585 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.740 0.770 7.660 1.000 ;
        RECT  4.355 0.885 5.970 1.115 ;
        RECT  7.375 0.770 7.660 1.600 ;
        RECT  2.125 3.420 2.410 3.760 ;
        RECT  4.450 3.385 6.330 3.615 ;
        RECT  2.125 3.530 3.580 3.760 ;
        RECT  7.520 3.365 7.860 3.845 ;
        RECT  6.100 3.615 7.860 3.845 ;
        RECT  4.450 3.385 4.680 3.885 ;
        RECT  3.365 3.655 4.680 3.885 ;
        RECT  9.335 0.780 10.485 1.010 ;
        RECT  8.020 0.630 8.360 1.430 ;
        RECT  9.335 0.780 9.565 1.430 ;
        RECT  7.890 1.200 9.565 1.430 ;
        RECT  6.780 1.885 8.120 2.115 ;
        RECT  6.780 1.800 7.065 2.180 ;
        RECT  10.255 0.780 10.485 2.770 ;
        RECT  7.890 1.200 8.120 3.005 ;
        RECT  10.255 2.460 11.375 2.770 ;
        RECT  7.890 2.665 8.360 3.005 ;
        RECT  11.190 1.795 11.840 2.135 ;
        RECT  8.350 2.020 8.715 2.360 ;
        RECT  8.525 2.225 8.820 2.440 ;
        RECT  8.590 2.225 8.820 2.910 ;
        RECT  11.610 1.795 11.840 3.230 ;
        RECT  8.590 2.680 10.025 2.910 ;
        RECT  9.795 1.240 10.025 3.230 ;
        RECT  11.610 2.890 12.050 3.230 ;
        RECT  9.795 3.000 12.050 3.230 ;
        RECT  10.715 0.630 13.040 0.860 ;
        RECT  10.715 0.630 11.000 1.005 ;
        RECT  12.700 0.630 13.040 1.195 ;
        RECT  11.470 1.090 12.300 1.430 ;
        RECT  12.070 1.090 12.300 2.385 ;
        RECT  12.280 2.155 12.515 3.145 ;
        RECT  13.760 2.740 14.045 3.090 ;
        RECT  12.280 2.860 14.045 3.090 ;
        RECT  12.280 2.860 13.580 3.145 ;
        RECT  12.280 2.155 12.510 3.750 ;
        RECT  11.320 3.460 12.510 3.750 ;
        RECT  12.530 1.495 12.815 1.835 ;
        RECT  12.530 1.605 14.400 1.835 ;
        RECT  14.060 1.660 14.510 1.945 ;
        RECT  14.275 1.660 14.510 2.640 ;
        RECT  14.275 2.300 14.775 2.640 ;
        RECT  14.275 1.660 14.505 3.550 ;
        RECT  13.820 3.320 14.505 3.550 ;
        RECT  13.820 3.320 14.050 4.160 ;
        RECT  13.710 3.820 14.050 4.160 ;
        RECT  1.255 1.585 2.40 1.815 ;
        RECT  4.450 2.870 5.90 3.155 ;
        RECT  4.450 2.925 6.30 3.155 ;
        RECT  2.255 0.630 3.20 0.860 ;
        RECT  9.795 3.000 11.80 3.230 ;
        RECT  10.715 0.630 12.60 0.860 ;
    END
END SDFFRX1

MACRO SDFFRX0
    CLASS CORE ;
    FOREIGN SDFFRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.225 1.260 15.625 4.150 ;
        RECT  15.100 1.260 15.625 1.600 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.550  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.300 2.860 14.995 3.350 ;
        RECT  14.765 1.830 14.995 3.350 ;
        RECT  14.515 1.830 14.995 2.060 ;
        RECT  14.515 0.630 14.745 2.060 ;
        RECT  14.200 0.630 14.745 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.302  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.245 13.225 2.820 ;
        END
    END RN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.830 2.215 9.325 2.720 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  14.300 3.810 14.680 5.280 ;
        RECT  12.235 3.910 12.570 5.280 ;
        RECT  9.510 3.630 9.850 5.280 ;
        RECT  8.310 3.910 8.650 5.280 ;
        RECT  4.830 3.865 5.170 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.100 -0.400 15.440 0.800 ;
        RECT  13.400 -0.400 13.740 0.950 ;
        RECT  8.615 -0.400 8.900 1.515 ;
        RECT  4.485 -0.400 4.825 0.655 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.815 ;
        RECT  2.930 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  3.500 1.345 5.425 1.575 ;
        RECT  3.505 1.805 5.520 2.090 ;
        RECT  5.235 1.805 5.520 2.180 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.750 1.230 6.655 1.540 ;
        RECT  3.965 2.325 4.950 2.665 ;
        RECT  4.605 2.325 4.950 3.175 ;
        RECT  4.605 2.945 5.980 3.175 ;
        RECT  5.750 1.230 5.980 3.175 ;
        RECT  5.805 3.025 6.500 3.255 ;
        RECT  6.270 3.025 6.500 3.790 ;
        RECT  6.270 3.450 6.610 3.790 ;
        RECT  4.370 3.405 5.610 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.420 3.440 5.650 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.030 3.640 7.370 4.250 ;
        RECT  5.420 4.020 7.370 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  3.960 0.630 4.190 1.115 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  5.290 0.770 7.455 1.000 ;
        RECT  3.960 0.885 5.520 1.115 ;
        RECT  7.115 0.770 7.455 1.570 ;
        RECT  6.210 1.840 6.495 2.210 ;
        RECT  6.210 1.870 7.585 2.210 ;
        RECT  9.130 0.770 10.280 1.000 ;
        RECT  7.815 1.230 8.155 1.985 ;
        RECT  9.130 0.770 9.360 1.985 ;
        RECT  7.815 1.755 9.360 1.985 ;
        RECT  10.050 0.770 10.280 2.755 ;
        RECT  6.210 2.510 6.545 2.795 ;
        RECT  10.050 2.415 10.800 2.755 ;
        RECT  6.210 2.550 7.080 2.795 ;
        RECT  6.850 2.550 7.080 3.220 ;
        RECT  7.815 1.230 8.045 3.220 ;
        RECT  6.850 2.875 8.045 3.220 ;
        RECT  9.590 1.230 9.820 3.220 ;
        RECT  11.160 1.765 11.545 3.220 ;
        RECT  8.910 2.990 11.545 3.220 ;
        RECT  8.910 2.990 9.250 3.395 ;
        RECT  8.910 2.990 9.140 3.680 ;
        RECT  7.790 3.450 9.140 3.680 ;
        RECT  7.790 3.450 8.075 3.880 ;
        RECT  10.510 0.635 12.860 0.865 ;
        RECT  12.520 0.635 12.860 0.970 ;
        RECT  10.510 0.635 10.850 0.975 ;
        RECT  11.485 1.175 12.005 1.515 ;
        RECT  11.775 3.125 13.610 3.465 ;
        RECT  11.775 1.175 12.005 3.970 ;
        RECT  10.805 3.630 12.005 3.970 ;
        RECT  13.840 1.410 14.285 1.750 ;
        RECT  12.450 1.695 14.070 2.015 ;
        RECT  13.840 2.290 14.535 2.630 ;
        RECT  13.840 1.410 14.070 4.175 ;
        RECT  13.195 3.835 14.070 4.175 ;
        RECT  0.980 1.585 2.30 1.815 ;
        RECT  1.445 1.125 2.20 1.355 ;
        RECT  3.505 1.805 4.50 2.090 ;
        RECT  1.995 3.710 3.00 3.940 ;
        RECT  1.980 0.630 3.40 0.860 ;
        RECT  5.290 0.770 6.60 1.000 ;
        RECT  8.910 2.990 10.50 3.220 ;
        RECT  10.510 0.635 11.10 0.865 ;
    END
END SDFFRX0

MACRO SDFFRSX4
    CLASS CORE ;
    FOREIGN SDFFRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.680 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.105  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  22.160 1.130 22.500 3.295 ;
        RECT  20.830 2.250 22.500 2.630 ;
        RECT  20.830 2.250 21.205 3.295 ;
        RECT  20.830 1.130 21.060 3.295 ;
        RECT  20.720 1.130 21.060 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.135  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.155 3.010 20.585 3.240 ;
        RECT  20.355 1.700 20.585 3.240 ;
        RECT  18.055 1.700 20.585 1.930 ;
        RECT  19.595 3.010 19.935 3.350 ;
        RECT  19.280 1.130 19.620 1.930 ;
        RECT  18.155 2.860 18.775 3.240 ;
        RECT  18.155 2.860 18.495 4.030 ;
        RECT  18.055 1.130 18.285 1.930 ;
        RECT  17.840 1.130 18.285 1.470 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.225 1.640 16.885 2.020 ;
        RECT  16.225 1.640 16.565 2.130 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.185 2.190 15.685 2.690 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.955 1.645 10.585 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 22.680 0.400 ;
        RECT  21.440 -0.400 21.780 1.470 ;
        RECT  20.000 -0.400 20.340 1.470 ;
        RECT  18.560 -0.400 18.900 1.470 ;
        RECT  15.945 -0.400 16.285 0.950 ;
        RECT  10.350 -0.400 10.690 0.955 ;
        RECT  4.775 -0.400 6.345 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 22.680 5.280 ;
        RECT  21.520 3.530 21.860 5.280 ;
        RECT  20.225 3.685 20.565 5.280 ;
        RECT  18.875 3.470 19.215 5.280 ;
        RECT  17.395 4.070 17.735 5.280 ;
        RECT  14.955 3.910 16.415 5.280 ;
        RECT  12.655 3.965 12.995 5.280 ;
        RECT  10.235 2.910 10.535 5.280 ;
        RECT  4.830 3.965 6.300 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 6.485 2.095 ;
        RECT  6.255 1.860 6.485 2.800 ;
        RECT  6.255 2.460 6.595 2.800 ;
        RECT  3.895 1.815 4.125 3.370 ;
        RECT  3.895 3.085 4.260 3.370 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 7.055 1.585 ;
        RECT  5.445 1.355 7.055 1.630 ;
        RECT  6.765 1.355 7.055 1.695 ;
        RECT  7.285 1.160 8.330 1.500 ;
        RECT  4.355 2.325 5.600 2.665 ;
        RECT  5.260 2.325 5.600 3.275 ;
        RECT  7.285 1.160 7.515 3.540 ;
        RECT  5.260 3.045 7.515 3.275 ;
        RECT  7.200 3.200 7.545 3.540 ;
        RECT  4.450 3.505 6.820 3.735 ;
        RECT  6.590 3.505 6.820 4.000 ;
        RECT  2.020 3.600 4.640 3.830 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  8.010 2.980 8.350 4.000 ;
        RECT  6.590 3.770 8.350 4.000 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.640 0.700 8.790 0.930 ;
        RECT  4.315 0.895 6.870 1.125 ;
        RECT  8.560 0.700 8.790 1.660 ;
        RECT  8.560 1.320 9.145 1.660 ;
        RECT  10.920 0.775 12.070 1.005 ;
        RECT  9.020 0.735 9.890 1.090 ;
        RECT  9.385 0.735 9.890 1.415 ;
        RECT  10.920 0.775 11.150 1.415 ;
        RECT  9.385 1.185 11.150 1.415 ;
        RECT  11.840 0.775 12.070 2.090 ;
        RECT  11.840 1.860 13.505 2.090 ;
        RECT  10.815 1.185 11.135 2.100 ;
        RECT  9.385 0.735 9.615 2.150 ;
        RECT  13.165 1.860 13.505 2.200 ;
        RECT  9.260 1.920 9.545 3.195 ;
        RECT  7.745 1.800 8.055 2.160 ;
        RECT  7.745 1.890 9.030 2.160 ;
        RECT  11.380 1.240 11.610 2.680 ;
        RECT  11.380 2.340 12.025 2.680 ;
        RECT  13.835 1.670 14.135 2.680 ;
        RECT  9.775 2.450 14.135 2.680 ;
        RECT  10.915 2.450 11.255 2.860 ;
        RECT  8.690 1.890 9.030 3.655 ;
        RECT  10.915 2.450 11.145 3.855 ;
        RECT  9.775 2.450 10.005 3.655 ;
        RECT  8.690 3.425 10.005 3.655 ;
        RECT  12.125 3.505 13.635 3.735 ;
        RECT  13.405 3.505 13.635 4.100 ;
        RECT  10.915 3.625 12.355 3.855 ;
        RECT  13.405 3.760 13.745 4.100 ;
        RECT  12.300 0.630 15.485 0.860 ;
        RECT  14.675 0.630 15.485 0.950 ;
        RECT  12.300 0.630 12.595 1.500 ;
        RECT  13.420 1.100 13.760 1.440 ;
        RECT  13.420 1.210 14.595 1.440 ;
        RECT  17.025 2.270 17.365 2.610 ;
        RECT  16.375 2.380 17.365 2.610 ;
        RECT  14.365 1.210 14.595 3.275 ;
        RECT  16.375 2.380 16.605 3.275 ;
        RECT  11.465 3.045 16.605 3.275 ;
        RECT  15.515 3.045 15.855 3.385 ;
        RECT  11.465 3.045 11.805 3.395 ;
        RECT  13.975 3.045 14.265 3.780 ;
        RECT  14.825 1.180 17.480 1.410 ;
        RECT  14.825 1.180 15.165 1.675 ;
        RECT  17.140 1.180 17.480 2.040 ;
        RECT  17.140 1.810 17.825 2.040 ;
        RECT  17.595 2.250 20.125 2.480 ;
        RECT  19.785 2.250 20.125 2.590 ;
        RECT  17.595 1.810 17.825 3.070 ;
        RECT  16.835 2.840 17.825 3.070 ;
        RECT  16.835 2.840 17.175 3.660 ;
        RECT  1.145 1.585 2.40 1.815 ;
        RECT  3.895 1.860 5.60 2.095 ;
        RECT  1.605 1.125 3.40 1.355 ;
        RECT  3.855 1.355 6.80 1.585 ;
        RECT  5.260 3.045 6.40 3.275 ;
        RECT  4.450 3.505 5.40 3.735 ;
        RECT  2.020 3.600 3.30 3.830 ;
        RECT  2.255 0.630 3.20 0.895 ;
        RECT  6.640 0.700 7.80 0.930 ;
        RECT  4.315 0.895 5.80 1.125 ;
        RECT  9.775 2.450 13.80 2.680 ;
        RECT  12.300 0.630 14.30 0.860 ;
        RECT  11.465 3.045 15.70 3.275 ;
        RECT  14.825 1.180 16.30 1.410 ;
        RECT  17.595 2.250 19.70 2.480 ;
    END
END SDFFRSX4

MACRO SDFFRSX2
    CLASS CORE ;
    FOREIGN SDFFRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.650 0.820 16.885 3.240 ;
        RECT  16.340 2.860 16.735 4.180 ;
        RECT  16.500 0.820 16.885 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 2.035 14.125 2.375 ;
        RECT  13.355 2.035 13.735 2.630 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.050 14.995 2.630 ;
        RECT  14.475 2.050 14.995 2.395 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.765 1.230 18.160 2.020 ;
        RECT  17.660 2.640 18.000 3.550 ;
        RECT  17.765 1.230 18.000 3.550 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.995 2.020 9.370 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  18.380 -0.400 18.720 0.710 ;
        RECT  17.260 -0.400 17.600 0.710 ;
        RECT  15.740 -0.400 16.080 0.970 ;
        RECT  14.395 -0.400 14.735 0.890 ;
        RECT  9.385 -0.400 9.670 1.330 ;
        RECT  5.630 -0.400 5.920 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  18.380 2.640 18.720 5.280 ;
        RECT  17.100 3.950 17.440 5.280 ;
        RECT  15.580 4.170 15.920 5.280 ;
        RECT  14.260 3.910 14.600 5.280 ;
        RECT  13.120 3.825 13.460 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.965 3.900 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.265 1.630 ;
        RECT  4.135 1.550 4.475 2.090 ;
        RECT  3.895 1.860 6.545 2.090 ;
        RECT  6.205 1.860 6.545 2.375 ;
        RECT  3.895 1.860 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.850 1.190 7.495 1.530 ;
        RECT  4.355 2.320 5.645 2.635 ;
        RECT  6.850 1.190 7.080 3.210 ;
        RECT  5.305 2.320 5.645 3.210 ;
        RECT  6.850 2.870 7.475 3.210 ;
        RECT  5.305 2.980 7.475 3.210 ;
        RECT  4.505 3.440 6.705 3.670 ;
        RECT  2.120 3.500 4.735 3.730 ;
        RECT  7.895 3.535 8.235 3.845 ;
        RECT  6.475 3.615 8.235 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.150 0.725 8.295 0.955 ;
        RECT  5.170 0.940 6.380 1.170 ;
        RECT  7.955 0.725 8.295 1.600 ;
        RECT  9.900 0.800 11.050 1.030 ;
        RECT  8.610 0.630 8.950 1.790 ;
        RECT  10.820 0.800 11.050 1.790 ;
        RECT  9.900 0.800 10.130 1.790 ;
        RECT  8.535 1.560 10.130 1.790 ;
        RECT  10.820 1.560 12.475 1.790 ;
        RECT  12.135 1.560 12.475 1.895 ;
        RECT  8.535 1.560 8.765 2.845 ;
        RECT  8.240 2.020 8.765 2.360 ;
        RECT  9.700 1.560 10.040 2.360 ;
        RECT  8.425 2.020 8.765 2.845 ;
        RECT  7.310 1.800 7.650 2.115 ;
        RECT  7.310 1.885 7.970 2.115 ;
        RECT  11.245 2.120 11.585 2.460 ;
        RECT  11.245 2.225 12.630 2.460 ;
        RECT  10.360 2.230 12.630 2.460 ;
        RECT  12.345 2.225 12.630 2.565 ;
        RECT  7.740 1.885 7.970 3.305 ;
        RECT  9.030 2.860 10.590 3.145 ;
        RECT  10.360 1.260 10.590 3.145 ;
        RECT  7.740 3.075 9.260 3.305 ;
        RECT  11.280 0.630 13.975 0.860 ;
        RECT  13.635 0.630 13.975 1.105 ;
        RECT  11.280 0.630 11.565 1.330 ;
        RECT  12.405 1.090 13.090 1.330 ;
        RECT  12.860 1.090 13.090 3.090 ;
        RECT  13.965 2.605 14.305 3.090 ;
        RECT  15.225 2.750 15.565 3.090 ;
        RECT  11.725 2.860 15.565 3.090 ;
        RECT  11.725 2.860 12.065 3.615 ;
        RECT  13.355 1.380 13.705 1.720 ;
        RECT  13.355 1.490 15.765 1.720 ;
        RECT  15.425 1.490 15.765 2.210 ;
        RECT  15.425 1.870 16.285 2.210 ;
        RECT  15.795 1.870 16.025 3.720 ;
        RECT  15.020 3.380 16.025 3.720 ;
        RECT  1.255 1.585 2.10 1.815 ;
        RECT  2.825 1.090 3.30 1.320 ;
        RECT  1.715 1.125 2.20 1.355 ;
        RECT  3.895 1.860 5.80 2.090 ;
        RECT  5.305 2.980 6.60 3.210 ;
        RECT  4.505 3.440 5.60 3.670 ;
        RECT  2.120 3.500 3.90 3.730 ;
        RECT  2.255 0.630 4.80 0.860 ;
        RECT  6.150 0.725 7.20 0.955 ;
        RECT  10.360 2.230 11.80 2.460 ;
        RECT  11.280 0.630 12.30 0.860 ;
        RECT  11.725 2.860 14.70 3.090 ;
        RECT  13.355 1.490 14.30 1.720 ;
    END
END SDFFRSX2

MACRO SDFFRSX1
    CLASS CORE ;
    FOREIGN SDFFRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 2.860 17.515 3.240 ;
        RECT  17.120 0.940 17.460 1.280 ;
        RECT  17.120 2.860 17.450 4.180 ;
        RECT  17.120 0.940 17.350 4.180 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.425 1.640 16.885 2.020 ;
        RECT  15.885 2.870 16.655 3.100 ;
        RECT  16.425 1.235 16.655 3.100 ;
        RECT  15.840 1.235 16.655 1.465 ;
        RECT  15.670 3.680 16.115 3.965 ;
        RECT  15.885 2.870 16.115 3.965 ;
        RECT  15.840 0.700 16.070 1.465 ;
        RECT  15.700 3.660 16.115 3.965 ;
        RECT  15.680 0.700 16.070 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.665 3.995 2.030 4.250 ;
        RECT  1.665 3.960 2.010 4.250 ;
        RECT  1.665 3.470 1.895 4.250 ;
        RECT  1.410 3.470 1.895 3.815 ;
        RECT  1.385 3.470 1.895 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.970 2.800 3.655 3.190 ;
        RECT  2.970 2.045 3.200 3.190 ;
        RECT  0.575 2.045 3.200 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.805 2.650 3.190 ;
        RECT  2.310 2.580 2.650 3.190 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.310 2.045 14.040 2.580 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.460 1.930 15.090 2.580 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.995 2.020 9.400 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.005 ;
        RECT  14.385 -0.400 14.725 1.025 ;
        RECT  9.450 -0.400 9.755 0.970 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.390 3.330 16.730 5.280 ;
        RECT  15.085 4.170 15.425 5.280 ;
        RECT  13.295 3.665 13.635 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.855 3.845 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.720 1.815 ;
        RECT  3.380 1.555 3.720 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.310 1.630 ;
        RECT  4.140 1.550 4.480 2.090 ;
        RECT  3.950 1.860 6.710 2.090 ;
        RECT  6.370 1.860 6.710 2.460 ;
        RECT  3.950 1.860 4.180 3.135 ;
        RECT  3.930 2.795 4.270 3.135 ;
        RECT  6.955 1.200 7.540 1.540 ;
        RECT  4.420 2.320 5.535 2.605 ;
        RECT  5.305 2.320 5.535 3.155 ;
        RECT  6.955 1.200 7.185 3.385 ;
        RECT  5.305 2.870 7.185 3.155 ;
        RECT  6.955 3.045 7.510 3.385 ;
        RECT  4.380 3.385 6.725 3.615 ;
        RECT  2.125 3.420 4.505 3.650 ;
        RECT  2.125 3.420 2.410 3.760 ;
        RECT  7.930 3.535 8.270 3.845 ;
        RECT  6.495 3.615 8.270 3.845 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.740 8.230 0.970 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  8.000 0.740 8.230 1.600 ;
        RECT  8.000 1.260 8.305 1.600 ;
        RECT  7.415 1.800 7.700 2.700 ;
        RECT  7.415 2.470 7.970 2.700 ;
        RECT  10.445 1.240 10.675 3.120 ;
        RECT  9.990 2.625 10.675 3.120 ;
        RECT  7.740 2.470 7.970 3.305 ;
        RECT  9.115 2.890 11.785 3.120 ;
        RECT  11.445 2.890 11.785 3.230 ;
        RECT  7.740 3.075 9.345 3.305 ;
        RECT  9.985 0.780 11.135 1.010 ;
        RECT  8.650 0.630 8.990 1.430 ;
        RECT  8.650 1.200 10.215 1.430 ;
        RECT  9.985 0.780 10.215 1.430 ;
        RECT  8.535 1.205 8.765 2.845 ;
        RECT  9.750 1.200 10.105 2.105 ;
        RECT  10.905 0.780 11.135 2.450 ;
        RECT  8.150 1.950 8.765 2.290 ;
        RECT  10.905 2.220 11.655 2.450 ;
        RECT  11.315 2.330 12.420 2.560 ;
        RECT  8.425 1.950 8.765 2.845 ;
        RECT  12.135 2.330 12.420 3.450 ;
        RECT  11.365 0.630 13.960 0.860 ;
        RECT  11.365 0.630 11.650 1.005 ;
        RECT  13.620 0.630 13.960 1.200 ;
        RECT  12.320 1.090 12.880 1.400 ;
        RECT  12.650 2.810 15.145 3.040 ;
        RECT  12.650 2.810 14.170 3.070 ;
        RECT  12.650 1.090 12.880 3.970 ;
        RECT  11.725 3.680 12.880 3.970 ;
        RECT  13.270 1.425 13.570 1.740 ;
        RECT  13.270 1.435 15.605 1.665 ;
        RECT  13.270 1.435 13.610 1.740 ;
        RECT  15.375 1.695 15.920 1.980 ;
        RECT  15.375 2.300 16.170 2.640 ;
        RECT  15.375 1.435 15.605 3.450 ;
        RECT  14.285 3.270 15.525 3.500 ;
        RECT  14.285 3.270 14.625 4.005 ;
        RECT  1.255 1.585 2.70 1.815 ;
        RECT  2.825 1.090 3.90 1.320 ;
        RECT  3.950 1.860 5.70 2.090 ;
        RECT  4.380 3.385 5.80 3.615 ;
        RECT  2.125 3.420 3.30 3.650 ;
        RECT  2.255 0.630 4.20 0.860 ;
        RECT  6.145 0.740 7.80 0.970 ;
        RECT  9.115 2.890 10.60 3.120 ;
        RECT  11.365 0.630 12.40 0.860 ;
        RECT  12.650 2.810 14.90 3.040 ;
        RECT  13.270 1.435 14.40 1.665 ;
    END
END SDFFRSX1

MACRO SDFFRSX0
    CLASS CORE ;
    FOREIGN SDFFRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.485 2.860 16.885 3.350 ;
        RECT  16.485 1.170 16.715 3.350 ;
        RECT  16.305 3.010 16.645 4.150 ;
        RECT  16.265 1.170 16.715 1.500 ;
        RECT  16.255 1.170 16.715 1.455 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.455  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.395 2.550 16.070 2.780 ;
        RECT  15.840 1.625 16.070 2.780 ;
        RECT  15.770 0.630 16.000 1.810 ;
        RECT  15.175 0.630 16.000 0.950 ;
        RECT  15.250 2.860 15.625 3.350 ;
        RECT  15.395 2.550 15.625 3.350 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.245 13.350 2.750 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 2.250 14.560 2.680 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.760 2.250 9.275 2.630 ;
        RECT  8.760 2.160 9.110 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.250 3.810 15.605 5.280 ;
        RECT  12.715 3.910 13.520 5.280 ;
        RECT  9.940 3.630 10.280 5.280 ;
        RECT  8.655 3.940 8.995 5.280 ;
        RECT  4.830 3.865 5.620 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.255 -0.400 16.595 0.710 ;
        RECT  14.145 -0.400 14.485 0.950 ;
        RECT  9.045 -0.400 9.330 1.400 ;
        RECT  4.715 -0.400 5.055 0.710 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.500 1.090 3.730 1.630 ;
        RECT  5.565 1.395 5.855 1.630 ;
        RECT  3.500 1.400 5.855 1.630 ;
        RECT  3.505 1.860 5.950 2.120 ;
        RECT  5.665 1.860 5.950 2.205 ;
        RECT  3.505 1.860 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  6.180 1.230 7.085 1.540 ;
        RECT  3.965 2.350 5.275 2.665 ;
        RECT  4.930 2.350 5.275 3.175 ;
        RECT  4.930 2.945 6.410 3.175 ;
        RECT  6.180 1.230 6.410 3.175 ;
        RECT  6.235 3.025 6.825 3.255 ;
        RECT  6.595 3.025 6.825 3.790 ;
        RECT  6.595 3.450 6.935 3.790 ;
        RECT  4.370 3.405 6.055 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.850 3.430 6.080 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.355 3.940 7.695 4.250 ;
        RECT  5.850 4.020 7.695 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  3.960 0.630 4.190 1.170 ;
        RECT  5.285 0.770 7.885 1.000 ;
        RECT  3.960 0.940 5.515 1.170 ;
        RECT  7.545 0.770 7.885 1.570 ;
        RECT  6.640 2.510 7.395 2.795 ;
        RECT  10.020 1.230 10.250 3.360 ;
        RECT  10.020 3.020 11.230 3.360 ;
        RECT  8.425 3.110 11.230 3.360 ;
        RECT  8.425 3.110 9.595 3.450 ;
        RECT  7.165 2.510 7.395 3.710 ;
        RECT  8.425 3.110 8.655 3.710 ;
        RECT  7.165 3.480 8.655 3.710 ;
        RECT  9.560 0.770 10.710 1.000 ;
        RECT  8.245 1.230 8.585 1.870 ;
        RECT  8.245 1.640 9.790 1.870 ;
        RECT  6.640 1.840 6.925 2.180 ;
        RECT  7.695 1.870 8.475 2.180 ;
        RECT  10.480 0.770 10.710 2.290 ;
        RECT  9.560 0.770 9.790 2.160 ;
        RECT  9.490 1.640 9.790 2.160 ;
        RECT  6.640 1.895 8.475 2.180 ;
        RECT  10.480 2.060 11.245 2.290 ;
        RECT  10.905 2.170 11.915 2.400 ;
        RECT  7.845 1.870 8.075 3.250 ;
        RECT  11.685 2.170 11.915 3.440 ;
        RECT  7.845 2.965 8.195 3.250 ;
        RECT  11.685 3.100 12.025 3.440 ;
        RECT  10.940 0.630 13.685 0.860 ;
        RECT  0.980 1.585 2.60 1.960 ;
        RECT  1.445 1.125 2.50 1.355 ;
        RECT  3.500 1.400 4.30 1.630 ;
        RECT  3.505 1.860 4.40 2.120 ;
        RECT  1.995 3.710 3.60 3.940 ;
        RECT  1.980 0.630 3.50 0.860 ;
        RECT  5.285 0.770 6.20 1.000 ;
        RECT  8.425 3.110 10.60 3.360 ;
        RECT  10.940 0.630 12.40 0.860 ;
        RECT  13.345 0.630 13.685 1.200 ;
        RECT  10.940 0.630 11.225 1.400 ;
        RECT  12.115 1.090 12.485 1.400 ;
        RECT  12.255 3.125 14.525 3.465 ;
        RECT  12.255 1.090 12.485 3.970 ;
        RECT  11.235 3.670 12.485 3.970 ;
        RECT  13.075 1.430 15.515 1.775 ;
        RECT  15.175 1.350 15.515 2.320 ;
        RECT  14.790 1.430 15.515 2.320 ;
        RECT  14.790 1.980 15.610 2.320 ;
        RECT  14.790 1.430 15.020 4.175 ;
        RECT  14.205 3.835 15.020 4.175 ;
    END
END SDFFRSX0

MACRO SDFFRSQX4
    CLASS CORE ;
    FOREIGN SDFFRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 1.130 19.980 4.030 ;
        RECT  18.200 2.250 19.980 2.630 ;
        RECT  18.200 1.130 18.540 4.030 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.875 1.640 16.365 2.150 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.175 2.180 15.645 2.700 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.005 1.640 10.535 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.470 ;
        RECT  17.440 -0.400 17.780 0.800 ;
        RECT  15.875 -0.400 16.215 0.760 ;
        RECT  10.305 -0.400 10.645 0.950 ;
        RECT  4.775 -0.400 6.345 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  18.920 2.860 19.260 5.280 ;
        RECT  17.440 4.070 17.780 5.280 ;
        RECT  14.955 3.910 16.415 5.280 ;
        RECT  12.655 3.965 12.995 5.280 ;
        RECT  10.235 2.910 10.535 5.280 ;
        RECT  4.830 3.965 6.300 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 6.485 2.095 ;
        RECT  6.255 1.860 6.485 2.800 ;
        RECT  6.255 2.460 6.595 2.800 ;
        RECT  3.895 1.815 4.125 3.370 ;
        RECT  3.895 3.085 4.260 3.370 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 7.055 1.585 ;
        RECT  5.445 1.355 7.055 1.630 ;
        RECT  6.765 1.355 7.055 1.695 ;
        RECT  7.285 1.160 8.285 1.500 ;
        RECT  4.355 2.325 4.640 2.665 ;
        RECT  4.355 2.435 5.490 2.665 ;
        RECT  5.260 2.435 5.490 3.275 ;
        RECT  5.260 2.935 5.600 3.275 ;
        RECT  7.285 1.160 7.515 3.540 ;
        RECT  5.260 3.045 7.515 3.275 ;
        RECT  7.200 3.200 7.545 3.540 ;
        RECT  4.450 3.505 6.820 3.735 ;
        RECT  6.590 3.505 6.820 4.000 ;
        RECT  2.020 3.600 4.640 3.830 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  8.010 2.980 8.350 4.000 ;
        RECT  6.590 3.770 8.350 4.000 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.640 0.700 8.745 0.930 ;
        RECT  4.315 0.895 6.870 1.125 ;
        RECT  8.515 0.700 8.745 1.660 ;
        RECT  8.515 1.320 9.145 1.660 ;
        RECT  10.875 0.775 12.025 1.005 ;
        RECT  8.975 0.735 9.845 1.090 ;
        RECT  9.375 0.735 9.845 1.410 ;
        RECT  9.375 1.180 11.105 1.410 ;
        RECT  11.795 0.775 12.025 2.090 ;
        RECT  11.795 1.860 13.450 2.090 ;
        RECT  10.875 0.775 11.105 2.100 ;
        RECT  10.765 1.180 11.105 2.100 ;
        RECT  9.375 0.735 9.605 2.150 ;
        RECT  13.110 1.860 13.450 2.200 ;
        RECT  9.260 1.920 9.545 3.195 ;
        RECT  7.745 1.890 9.000 2.120 ;
        RECT  7.745 1.765 8.055 2.160 ;
        RECT  11.335 1.240 11.565 2.680 ;
        RECT  11.335 2.340 12.025 2.680 ;
        RECT  13.790 1.670 14.075 2.680 ;
        RECT  9.775 2.450 14.075 2.680 ;
        RECT  10.915 2.450 11.255 2.860 ;
        RECT  8.700 1.890 9.000 3.655 ;
        RECT  10.915 2.450 11.145 3.855 ;
        RECT  9.775 2.450 10.005 3.655 ;
        RECT  8.700 3.425 10.005 3.655 ;
        RECT  12.125 3.505 13.635 3.735 ;
        RECT  13.405 3.505 13.635 4.100 ;
        RECT  10.915 3.625 12.355 3.855 ;
        RECT  13.405 3.760 13.745 4.100 ;
        RECT  12.255 0.630 15.210 0.860 ;
        RECT  14.870 0.630 15.210 0.950 ;
        RECT  12.255 0.630 12.550 1.500 ;
        RECT  13.360 1.100 13.700 1.440 ;
        RECT  13.360 1.210 14.535 1.440 ;
        RECT  17.025 2.270 17.365 2.610 ;
        RECT  16.375 2.380 17.365 2.610 ;
        RECT  14.305 1.210 14.535 3.275 ;
        RECT  16.375 2.380 16.605 3.275 ;
        RECT  11.465 3.045 16.605 3.275 ;
        RECT  15.515 3.045 15.855 3.385 ;
        RECT  11.465 3.045 11.805 3.395 ;
        RECT  13.975 3.045 14.265 3.780 ;
        RECT  14.765 1.180 17.280 1.410 ;
        RECT  16.940 1.350 17.825 1.580 ;
        RECT  14.765 1.180 15.095 1.730 ;
        RECT  17.595 1.350 17.825 3.070 ;
        RECT  16.835 2.840 17.825 3.070 ;
        RECT  16.835 2.840 17.175 3.660 ;
        RECT  1.145 1.585 2.80 1.815 ;
        RECT  3.895 1.860 5.80 2.095 ;
        RECT  1.605 1.125 3.70 1.355 ;
        RECT  3.855 1.355 6.00 1.585 ;
        RECT  5.260 3.045 6.60 3.275 ;
        RECT  4.450 3.505 5.50 3.735 ;
        RECT  2.020 3.600 3.60 3.830 ;
        RECT  2.255 0.630 3.60 0.895 ;
        RECT  6.640 0.700 7.30 0.930 ;
        RECT  4.315 0.895 5.20 1.125 ;
        RECT  9.775 2.450 13.40 2.680 ;
        RECT  12.255 0.630 14.80 0.860 ;
        RECT  11.465 3.045 15.40 3.275 ;
        RECT  14.765 1.180 16.90 1.410 ;
    END
END SDFFRSQX4

MACRO SDFFRSQX2
    CLASS CORE ;
    FOREIGN SDFFRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.560 1.240 16.900 2.630 ;
        RECT  16.340 2.250 16.735 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 2.035 14.125 2.375 ;
        RECT  13.355 2.035 13.735 2.630 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.050 14.995 2.630 ;
        RECT  14.475 2.050 14.995 2.395 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.995 2.020 9.370 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  17.120 -0.400 17.460 0.720 ;
        RECT  16.000 -0.400 16.340 0.720 ;
        RECT  14.395 -0.400 14.735 0.970 ;
        RECT  9.385 -0.400 9.670 1.330 ;
        RECT  5.630 -0.400 5.920 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  17.060 3.270 17.400 5.280 ;
        RECT  15.580 4.170 15.920 5.280 ;
        RECT  14.260 3.910 14.600 5.280 ;
        RECT  13.120 3.825 13.460 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.965 3.900 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.265 1.630 ;
        RECT  4.135 1.550 4.475 2.090 ;
        RECT  3.895 1.860 6.545 2.090 ;
        RECT  6.205 1.860 6.545 2.375 ;
        RECT  3.895 1.860 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.850 1.190 7.495 1.530 ;
        RECT  4.355 2.320 5.645 2.635 ;
        RECT  6.850 1.190 7.080 3.210 ;
        RECT  5.305 2.320 5.645 3.210 ;
        RECT  6.850 2.870 7.500 3.210 ;
        RECT  5.305 2.980 7.500 3.210 ;
        RECT  4.505 3.440 6.705 3.670 ;
        RECT  2.120 3.500 4.735 3.730 ;
        RECT  7.920 3.535 8.260 3.845 ;
        RECT  6.475 3.615 8.260 3.845 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.150 0.730 8.295 0.960 ;
        RECT  5.170 0.940 6.380 1.170 ;
        RECT  7.955 0.730 8.295 1.600 ;
        RECT  9.900 0.800 11.050 1.030 ;
        RECT  8.610 0.630 8.950 1.790 ;
        RECT  10.820 0.800 11.050 1.790 ;
        RECT  9.900 0.800 10.130 1.790 ;
        RECT  8.530 1.560 10.130 1.790 ;
        RECT  10.820 1.560 12.475 1.790 ;
        RECT  12.135 1.560 12.475 1.895 ;
        RECT  8.530 1.560 8.760 2.845 ;
        RECT  8.240 2.020 8.760 2.360 ;
        RECT  9.700 1.560 10.040 2.360 ;
        RECT  8.420 2.020 8.760 2.845 ;
        RECT  7.310 1.795 7.650 2.115 ;
        RECT  7.310 1.885 7.970 2.115 ;
        RECT  11.245 2.120 11.585 2.460 ;
        RECT  11.245 2.225 12.630 2.460 ;
        RECT  10.360 2.230 12.630 2.460 ;
        RECT  12.345 2.225 12.630 2.565 ;
        RECT  7.740 1.885 7.970 3.305 ;
        RECT  9.030 2.860 10.590 3.145 ;
        RECT  10.360 1.260 10.590 3.145 ;
        RECT  7.740 3.075 9.260 3.305 ;
        RECT  11.280 0.630 13.975 0.860 ;
        RECT  13.635 0.630 13.975 1.105 ;
        RECT  11.280 0.630 11.565 1.330 ;
        RECT  12.405 1.090 13.090 1.330 ;
        RECT  12.860 1.090 13.090 3.090 ;
        RECT  13.965 2.605 14.305 3.090 ;
        RECT  15.225 2.750 15.565 3.090 ;
        RECT  11.725 2.860 15.565 3.090 ;
        RECT  11.725 2.860 12.065 3.615 ;
        RECT  15.225 0.630 15.565 1.610 ;
        RECT  13.355 1.380 16.025 1.610 ;
        RECT  13.355 1.380 13.700 1.720 ;
        RECT  15.795 1.380 16.025 3.610 ;
        RECT  15.020 3.380 16.025 3.610 ;
        RECT  15.020 3.380 15.360 3.720 ;
        RECT  1.255 1.585 2.50 1.815 ;
        RECT  2.825 1.090 3.60 1.320 ;
        RECT  1.715 1.125 2.80 1.355 ;
        RECT  3.895 1.860 5.50 2.090 ;
        RECT  5.305 2.980 6.70 3.210 ;
        RECT  4.505 3.440 5.70 3.670 ;
        RECT  2.120 3.500 3.30 3.730 ;
        RECT  2.255 0.630 4.20 0.860 ;
        RECT  6.150 0.730 7.60 0.960 ;
        RECT  10.360 2.230 11.80 2.460 ;
        RECT  11.280 0.630 12.90 0.860 ;
        RECT  11.725 2.860 14.50 3.090 ;
        RECT  13.355 1.380 15.60 1.610 ;
    END
END SDFFRSQX2

MACRO SDFFRSQX1
    CLASS CORE ;
    FOREIGN SDFFRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.718  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.875 2.250 16.380 2.635 ;
        RECT  16.150 1.235 16.380 2.635 ;
        RECT  15.840 1.235 16.380 1.465 ;
        RECT  15.670 3.680 16.115 3.965 ;
        RECT  15.875 2.250 16.115 3.965 ;
        RECT  15.840 0.700 16.070 1.465 ;
        RECT  15.700 3.660 16.115 3.965 ;
        RECT  15.680 0.700 16.070 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.665 3.995 2.030 4.250 ;
        RECT  1.665 3.960 2.010 4.250 ;
        RECT  1.665 3.470 1.895 4.250 ;
        RECT  1.410 3.470 1.895 3.815 ;
        RECT  1.385 3.470 1.895 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.970 2.800 3.655 3.190 ;
        RECT  2.970 2.045 3.200 3.190 ;
        RECT  0.575 2.045 3.200 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.310 2.045 14.040 2.580 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.460 1.930 15.090 2.580 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.995 2.020 9.400 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.400 -0.400 16.740 1.005 ;
        RECT  14.385 -0.400 14.725 1.025 ;
        RECT  9.450 -0.400 9.755 0.970 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.390 3.330 16.730 5.280 ;
        RECT  15.085 4.170 15.425 5.280 ;
        RECT  13.295 3.665 13.635 5.280 ;
        RECT  10.530 3.480 10.870 5.280 ;
        RECT  9.230 3.535 9.570 5.280 ;
        RECT  4.855 3.845 6.245 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.720 1.815 ;
        RECT  3.380 1.555 3.720 1.895 ;
        RECT  0.115 1.240 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  4.710 1.090 4.940 1.630 ;
        RECT  4.710 1.400 6.310 1.630 ;
        RECT  4.140 1.550 4.480 2.090 ;
        RECT  3.950 1.860 6.710 2.090 ;
        RECT  6.370 1.860 6.710 2.460 ;
        RECT  3.950 1.860 4.180 3.135 ;
        RECT  3.930 2.795 4.270 3.135 ;
        RECT  6.955 1.200 7.540 1.540 ;
        RECT  4.420 2.320 5.535 2.605 ;
        RECT  5.305 2.320 5.535 3.155 ;
        RECT  6.955 1.200 7.185 3.385 ;
        RECT  5.305 2.870 7.185 3.155 ;
        RECT  6.955 3.045 7.510 3.385 ;
        RECT  4.380 3.385 6.725 3.615 ;
        RECT  2.125 3.420 4.505 3.650 ;
        RECT  2.125 3.420 2.410 3.760 ;
        RECT  7.930 3.535 8.270 3.845 ;
        RECT  6.495 3.615 8.270 3.845 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.740 8.305 0.970 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  8.000 0.740 8.305 1.600 ;
        RECT  7.415 1.820 7.700 2.700 ;
        RECT  7.415 2.470 7.970 2.700 ;
        RECT  9.990 2.715 10.675 3.120 ;
        RECT  10.445 1.240 10.675 3.120 ;
        RECT  9.115 2.865 10.675 3.120 ;
        RECT  7.740 2.470 7.970 3.305 ;
        RECT  9.115 2.890 11.785 3.120 ;
        RECT  11.445 2.890 11.785 3.230 ;
        RECT  7.740 3.075 9.345 3.305 ;
        RECT  9.985 0.780 11.135 1.010 ;
        RECT  8.650 0.630 8.990 1.430 ;
        RECT  9.985 0.780 10.215 1.430 ;
        RECT  8.535 1.200 10.215 1.430 ;
        RECT  8.535 1.200 8.765 2.845 ;
        RECT  9.750 1.200 10.105 2.120 ;
        RECT  10.905 0.780 11.135 2.450 ;
        RECT  8.150 1.950 8.765 2.290 ;
        RECT  10.905 2.220 11.655 2.450 ;
        RECT  11.315 2.330 12.420 2.560 ;
        RECT  8.425 1.950 8.765 2.845 ;
        RECT  12.135 2.330 12.420 3.450 ;
        RECT  11.365 0.630 13.960 0.860 ;
        RECT  11.365 0.630 11.650 1.005 ;
        RECT  13.620 0.630 13.960 1.200 ;
        RECT  12.320 1.090 12.880 1.400 ;
        RECT  12.650 2.810 15.145 3.040 ;
        RECT  12.650 2.810 14.170 3.070 ;
        RECT  12.650 1.090 12.880 3.970 ;
        RECT  11.725 3.680 12.880 3.970 ;
        RECT  13.270 1.425 13.570 1.740 ;
        RECT  13.270 1.435 15.605 1.665 ;
        RECT  13.270 1.435 13.610 1.740 ;
        RECT  15.375 1.695 15.920 1.980 ;
        RECT  15.375 1.435 15.605 3.450 ;
        RECT  14.285 3.270 15.525 3.500 ;
        RECT  14.285 3.270 14.625 4.005 ;
        RECT  1.255 1.585 2.70 1.815 ;
        RECT  2.825 1.090 3.60 1.320 ;
        RECT  3.950 1.860 5.90 2.090 ;
        RECT  4.380 3.385 5.70 3.615 ;
        RECT  2.125 3.420 3.60 3.650 ;
        RECT  2.255 0.630 4.70 0.860 ;
        RECT  6.145 0.740 7.60 0.970 ;
        RECT  9.115 2.890 10.80 3.120 ;
        RECT  11.365 0.630 12.30 0.860 ;
        RECT  12.650 2.810 14.40 3.040 ;
        RECT  13.270 1.435 14.60 1.665 ;
    END
END SDFFRSQX1

MACRO SDFFRSQX0
    CLASS CORE ;
    FOREIGN SDFFRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.512  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.220 2.860 15.635 3.350 ;
        RECT  15.405 0.635 15.635 3.350 ;
        RECT  14.855 0.635 15.635 0.975 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.590 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.286  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.245 13.380 2.895 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.985 2.250 14.485 2.795 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.760 2.250 9.275 2.630 ;
        RECT  8.760 2.160 9.110 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.220 3.810 15.560 5.280 ;
        RECT  12.715 3.910 13.520 5.280 ;
        RECT  9.940 3.630 10.280 5.280 ;
        RECT  8.655 3.940 8.995 5.280 ;
        RECT  4.830 3.865 5.620 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  13.825 -0.400 14.165 0.975 ;
        RECT  9.045 -0.400 9.330 1.400 ;
        RECT  4.715 -0.400 5.055 0.710 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.500 1.090 3.730 1.630 ;
        RECT  5.565 1.395 5.855 1.630 ;
        RECT  3.500 1.400 5.855 1.630 ;
        RECT  3.505 1.860 5.950 2.120 ;
        RECT  5.665 1.860 5.950 2.205 ;
        RECT  3.505 1.860 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  6.180 1.230 7.085 1.540 ;
        RECT  3.965 2.350 5.275 2.665 ;
        RECT  4.930 2.350 5.275 3.175 ;
        RECT  4.930 2.945 6.410 3.175 ;
        RECT  6.180 1.230 6.410 3.175 ;
        RECT  6.235 3.025 6.825 3.240 ;
        RECT  6.250 3.025 6.825 3.255 ;
        RECT  6.595 3.025 6.825 3.790 ;
        RECT  6.595 3.450 6.935 3.790 ;
        RECT  4.370 3.405 6.065 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.850 3.420 6.080 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.355 3.940 7.695 4.250 ;
        RECT  5.850 4.020 7.695 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  3.960 0.630 4.190 1.170 ;
        RECT  5.285 0.770 7.885 1.000 ;
        RECT  3.960 0.940 5.515 1.170 ;
        RECT  7.545 0.770 7.885 1.570 ;
        RECT  6.640 2.510 6.975 2.795 ;
        RECT  6.640 2.565 7.395 2.795 ;
        RECT  10.020 1.230 10.250 3.395 ;
        RECT  10.020 3.020 11.230 3.395 ;
        RECT  8.425 3.110 11.230 3.395 ;
        RECT  8.425 3.110 9.595 3.450 ;
        RECT  7.165 2.565 7.395 3.710 ;
        RECT  8.425 3.110 8.655 3.710 ;
        RECT  7.165 3.480 8.655 3.710 ;
        RECT  9.560 0.770 10.710 1.000 ;
        RECT  8.245 1.230 8.585 1.870 ;
        RECT  8.245 1.640 9.790 1.870 ;
        RECT  6.640 1.840 6.925 2.180 ;
        RECT  7.695 1.870 8.475 2.180 ;
        RECT  9.560 0.770 9.790 2.160 ;
        RECT  9.500 1.640 9.790 2.160 ;
        RECT  6.640 1.895 8.475 2.180 ;
        RECT  10.480 0.770 10.710 2.425 ;
        RECT  10.480 2.195 11.230 2.425 ;
        RECT  10.890 2.305 12.025 2.535 ;
        RECT  7.845 1.870 8.195 3.250 ;
        RECT  11.685 2.305 12.025 3.450 ;
        RECT  10.940 0.635 13.280 0.865 ;
        RECT  12.940 0.635 13.280 0.970 ;
        RECT  10.940 0.635 11.225 0.975 ;
        RECT  11.915 1.175 12.485 1.515 ;
        RECT  13.235 3.125 14.525 3.465 ;
        RECT  12.255 3.235 14.525 3.465 ;
        RECT  12.255 1.175 12.485 3.970 ;
        RECT  11.235 3.680 12.485 3.970 ;
        RECT  14.760 1.350 15.175 1.690 ;
        RECT  12.875 1.730 14.990 2.015 ;
        RECT  14.760 1.350 14.990 4.175 ;
        RECT  14.160 3.835 14.990 4.175 ;
        RECT  0.980 1.585 2.70 1.960 ;
        RECT  1.445 1.125 2.60 1.355 ;
        RECT  3.500 1.400 4.60 1.630 ;
        RECT  3.505 1.860 4.90 2.120 ;
        RECT  1.995 3.710 3.70 3.940 ;
        RECT  1.980 0.630 3.00 0.860 ;
        RECT  5.285 0.770 6.30 1.000 ;
        RECT  8.425 3.110 10.20 3.395 ;
        RECT  10.940 0.635 12.70 0.865 ;
        RECT  12.255 3.235 13.70 3.465 ;
        RECT  12.875 1.730 13.60 2.015 ;
    END
END SDFFRSQX0

MACRO SDFFRQX4
    CLASS CORE ;
    FOREIGN SDFFRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.010 1.130 19.350 4.010 ;
        RECT  17.570 2.250 19.350 2.630 ;
        RECT  17.570 1.130 17.910 4.010 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.020 1.640 15.625 2.100 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.505 1.660 9.965 2.160 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.290 -0.400 18.630 1.470 ;
        RECT  16.810 -0.400 17.150 0.725 ;
        RECT  15.500 -0.400 15.840 0.950 ;
        RECT  9.920 -0.400 10.205 0.970 ;
        RECT  4.775 -0.400 5.915 0.665 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.290 2.860 18.630 5.280 ;
        RECT  16.850 2.770 17.190 5.280 ;
        RECT  14.155 3.760 15.615 5.280 ;
        RECT  12.095 3.980 12.435 5.280 ;
        RECT  9.540 2.950 9.825 5.280 ;
        RECT  4.660 4.115 5.700 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.625 1.815 ;
        RECT  3.335 1.635 3.630 1.930 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.815 4.625 2.095 ;
        RECT  3.895 1.860 5.885 2.095 ;
        RECT  5.655 1.860 5.885 2.800 ;
        RECT  5.655 2.460 5.995 2.800 ;
        RECT  3.895 1.815 4.125 3.425 ;
        RECT  3.895 3.085 4.260 3.425 ;
        RECT  1.425 0.630 1.835 0.950 ;
        RECT  1.605 0.630 1.835 1.355 ;
        RECT  1.605 1.125 4.085 1.355 ;
        RECT  3.855 1.355 6.625 1.585 ;
        RECT  5.015 1.355 6.625 1.630 ;
        RECT  6.335 1.355 6.625 1.695 ;
        RECT  2.020 3.655 6.390 3.885 ;
        RECT  2.020 3.600 2.310 3.940 ;
        RECT  6.160 3.850 7.710 4.080 ;
        RECT  7.370 3.850 7.710 4.190 ;
        RECT  6.855 1.160 7.900 1.500 ;
        RECT  4.355 2.325 4.640 2.665 ;
        RECT  4.355 2.435 4.890 2.665 ;
        RECT  4.660 2.435 4.890 3.425 ;
        RECT  4.660 3.085 5.000 3.425 ;
        RECT  4.660 3.195 7.085 3.425 ;
        RECT  6.855 1.160 7.085 3.540 ;
        RECT  6.745 3.195 7.085 3.540 ;
        RECT  2.255 0.630 4.545 0.895 ;
        RECT  6.210 0.700 8.360 0.930 ;
        RECT  4.315 0.895 6.440 1.125 ;
        RECT  8.130 0.700 8.360 1.660 ;
        RECT  8.130 1.320 8.715 1.660 ;
        RECT  10.435 0.775 11.585 1.005 ;
        RECT  8.590 0.735 9.460 1.090 ;
        RECT  8.955 0.735 9.460 1.430 ;
        RECT  10.435 0.775 10.665 1.430 ;
        RECT  8.955 1.200 10.665 1.430 ;
        RECT  11.355 0.775 11.585 2.090 ;
        RECT  11.355 1.860 13.020 2.090 ;
        RECT  10.195 1.200 10.555 2.100 ;
        RECT  8.955 0.735 9.185 2.150 ;
        RECT  8.620 1.920 9.185 2.150 ;
        RECT  12.680 1.860 13.020 2.200 ;
        RECT  8.620 1.920 8.850 3.580 ;
        RECT  8.510 3.235 8.850 3.580 ;
        RECT  13.350 1.670 13.690 2.010 ;
        RECT  7.315 1.795 7.625 2.160 ;
        RECT  10.895 1.240 11.125 2.680 ;
        RECT  10.895 2.340 11.485 2.680 ;
        RECT  13.350 1.670 13.580 2.680 ;
        RECT  9.080 2.450 13.580 2.680 ;
        RECT  7.395 1.795 7.625 3.095 ;
        RECT  7.395 2.865 8.280 3.095 ;
        RECT  10.205 2.450 10.545 3.915 ;
        RECT  11.565 3.520 12.895 3.750 ;
        RECT  8.050 2.865 8.280 4.040 ;
        RECT  12.665 3.520 12.895 4.200 ;
        RECT  10.205 3.685 11.795 3.915 ;
        RECT  9.080 2.450 9.310 4.040 ;
        RECT  8.050 3.810 9.310 4.040 ;
        RECT  12.665 3.860 13.185 4.200 ;
        RECT  11.815 0.630 15.040 0.860 ;
        RECT  14.230 0.630 15.040 0.950 ;
        RECT  11.815 0.630 12.110 1.500 ;
        RECT  12.920 1.090 13.260 1.440 ;
        RECT  12.920 1.210 14.150 1.440 ;
        RECT  15.800 2.250 16.140 2.590 ;
        RECT  13.920 2.360 16.140 2.590 ;
        RECT  14.715 2.360 15.055 3.150 ;
        RECT  13.920 1.210 14.150 3.215 ;
        RECT  10.905 2.985 14.150 3.215 ;
        RECT  10.905 2.985 11.245 3.455 ;
        RECT  13.125 2.985 13.465 3.630 ;
        RECT  14.380 1.180 16.600 1.410 ;
        RECT  16.260 1.080 16.600 1.420 ;
        RECT  14.380 1.180 14.720 1.680 ;
        RECT  16.370 1.080 16.600 3.640 ;
        RECT  16.130 2.820 16.600 3.640 ;
        RECT  1.145 1.585 2.50 1.815 ;
        RECT  1.605 1.125 3.80 1.355 ;
        RECT  3.855 1.355 5.20 1.585 ;
        RECT  2.020 3.655 5.30 3.885 ;
        RECT  4.660 3.195 6.20 3.425 ;
        RECT  2.255 0.630 3.50 0.895 ;
        RECT  6.210 0.700 7.10 0.930 ;
        RECT  4.315 0.895 5.40 1.125 ;
        RECT  9.080 2.450 12.80 2.680 ;
        RECT  11.815 0.630 14.40 0.860 ;
        RECT  13.920 2.360 15.40 2.590 ;
        RECT  10.905 2.985 13.30 3.215 ;
        RECT  14.380 1.180 15.20 1.410 ;
    END
END SDFFRQX4

MACRO SDFFRQX2
    CLASS CORE ;
    FOREIGN SDFFRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.020 0.820 16.255 3.240 ;
        RECT  15.770 2.860 16.110 3.830 ;
        RECT  15.770 0.820 16.255 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.675 2.615 3.240 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        RECT  2.965 2.250 3.305 3.020 ;
        RECT  0.575 2.045 2.980 2.275 ;
        RECT  2.750 2.250 3.655 2.480 ;
        RECT  0.575 1.715 0.920 2.275 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.200 2.110 13.735 2.675 ;
        END
    END RN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.425 2.300 8.865 2.685 ;
        RECT  8.315 2.300 8.865 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 1.160 ;
        RECT  15.050 -0.400 15.390 1.160 ;
        RECT  14.005 -0.400 14.345 1.220 ;
        RECT  9.035 -0.400 9.320 1.330 ;
        RECT  5.630 -0.400 5.915 0.710 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.490 2.920 16.830 5.280 ;
        RECT  15.010 3.775 15.350 5.280 ;
        RECT  12.745 3.365 13.085 5.280 ;
        RECT  9.895 3.525 10.235 5.280 ;
        RECT  8.595 3.810 8.935 5.280 ;
        RECT  4.655 3.960 5.645 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.545 1.815 ;
        RECT  3.205 1.585 3.545 1.930 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.330 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  1.425 0.630 1.945 0.950 ;
        RECT  1.715 0.630 1.945 1.355 ;
        RECT  2.825 1.090 4.940 1.320 ;
        RECT  1.715 1.125 3.825 1.355 ;
        RECT  4.710 1.090 4.940 1.685 ;
        RECT  4.710 1.400 5.915 1.685 ;
        RECT  4.135 1.550 4.475 2.180 ;
        RECT  3.895 1.950 6.165 2.180 ;
        RECT  5.825 1.950 6.165 2.375 ;
        RECT  3.895 1.950 4.125 3.270 ;
        RECT  3.895 2.930 4.255 3.270 ;
        RECT  6.805 1.260 7.145 1.600 ;
        RECT  6.495 1.370 7.145 1.600 ;
        RECT  4.415 2.410 5.045 2.750 ;
        RECT  4.705 2.410 5.045 3.270 ;
        RECT  6.495 1.370 6.725 3.270 ;
        RECT  4.705 3.040 6.875 3.270 ;
        RECT  6.535 3.040 6.875 3.625 ;
        RECT  2.120 3.500 6.305 3.730 ;
        RECT  6.075 3.500 6.305 4.125 ;
        RECT  2.120 3.500 2.410 4.020 ;
        RECT  7.295 3.810 7.635 4.125 ;
        RECT  6.075 3.895 7.635 4.125 ;
        RECT  2.255 0.630 5.400 0.860 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.170 0.630 5.400 1.170 ;
        RECT  6.145 0.800 7.945 1.030 ;
        RECT  5.170 0.940 6.375 1.170 ;
        RECT  7.605 0.800 7.945 1.600 ;
        RECT  9.550 0.800 10.700 1.030 ;
        RECT  8.260 0.630 8.600 1.790 ;
        RECT  10.470 0.800 10.700 1.790 ;
        RECT  9.550 0.800 9.780 1.790 ;
        RECT  8.260 1.560 9.780 1.790 ;
        RECT  10.470 1.560 12.125 1.790 ;
        RECT  11.785 1.560 12.125 1.895 ;
        RECT  8.260 0.630 8.490 2.060 ;
        RECT  7.755 1.830 8.490 2.060 ;
        RECT  7.755 1.830 8.065 2.170 ;
        RECT  9.360 1.560 9.700 2.630 ;
        RECT  7.825 1.830 8.065 3.120 ;
        RECT  7.825 2.810 8.165 3.120 ;
        RECT  6.955 1.910 7.335 2.270 ;
        RECT  10.810 2.225 12.320 2.565 ;
        RECT  10.010 2.230 12.320 2.565 ;
        RECT  10.010 1.260 10.240 3.165 ;
        RECT  9.280 2.860 10.240 3.165 ;
        RECT  7.105 1.910 7.335 3.580 ;
        RECT  9.280 2.860 9.525 3.580 ;
        RECT  7.105 3.350 9.525 3.580 ;
        RECT  10.930 0.630 13.625 0.860 ;
        RECT  13.285 0.630 13.625 1.105 ;
        RECT  10.930 0.630 11.215 1.330 ;
        RECT  12.055 1.090 12.780 1.330 ;
        RECT  13.965 2.400 14.935 2.740 ;
        RECT  12.550 1.090 12.780 3.135 ;
        RECT  13.965 2.400 14.195 3.135 ;
        RECT  11.300 2.905 14.195 3.135 ;
        RECT  11.300 2.905 11.640 3.690 ;
        RECT  13.465 2.905 13.805 4.175 ;
        RECT  13.010 1.380 13.355 1.720 ;
        RECT  13.010 1.490 15.145 1.720 ;
        RECT  14.805 1.490 15.145 1.980 ;
        RECT  14.805 1.750 15.395 1.980 ;
        RECT  15.165 1.750 15.395 3.200 ;
        RECT  14.450 2.970 15.395 3.200 ;
        RECT  14.450 2.970 14.790 3.310 ;
        RECT  1.255 1.585 2.50 1.815 ;
        RECT  2.825 1.090 3.00 1.320 ;
        RECT  1.715 1.125 2.40 1.355 ;
        RECT  3.895 1.950 5.80 2.180 ;
        RECT  4.705 3.040 5.40 3.270 ;
        RECT  2.120 3.500 5.90 3.730 ;
        RECT  2.255 0.630 4.40 0.860 ;
        RECT  10.010 2.230 11.90 2.565 ;
        RECT  7.105 3.350 8.30 3.580 ;
        RECT  10.930 0.630 12.20 0.860 ;
        RECT  11.300 2.905 13.80 3.135 ;
        RECT  13.010 1.490 14.60 1.720 ;
    END
END SDFFRQX2

MACRO SDFFRQX1
    CLASS CORE ;
    FOREIGN SDFFRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.735 2.250 15.635 2.630 ;
        RECT  14.735 2.250 14.970 3.100 ;
        RECT  14.420 3.780 14.965 4.065 ;
        RECT  14.735 0.700 14.965 4.065 ;
        RECT  14.505 0.700 14.965 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 3.995 2.030 4.250 ;
        RECT  1.610 3.980 2.000 4.250 ;
        RECT  1.610 3.470 1.840 4.250 ;
        RECT  1.410 3.470 1.840 3.815 ;
        RECT  1.385 3.470 1.840 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.980 2.800 3.655 3.240 ;
        RECT  2.980 2.045 3.210 3.240 ;
        RECT  0.575 2.045 3.210 2.275 ;
        RECT  0.575 1.660 0.860 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.745 2.170 13.290 2.630 ;
        END
    END RN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.305 1.660 8.715 2.320 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  15.195 3.330 15.535 5.280 ;
        RECT  12.740 3.820 13.085 5.280 ;
        RECT  10.125 3.480 10.465 5.280 ;
        RECT  8.825 3.535 9.165 5.280 ;
        RECT  4.910 3.845 5.870 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.225 -0.400 15.565 1.040 ;
        RECT  13.470 -0.400 13.810 1.015 ;
        RECT  8.820 -0.400 9.105 0.970 ;
        RECT  4.815 -0.400 5.155 0.655 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.130 0.900 1.430 ;
        RECT  0.115 1.185 1.485 1.430 ;
        RECT  1.255 1.185 1.485 1.815 ;
        RECT  1.255 1.585 3.665 1.815 ;
        RECT  3.380 1.555 3.665 1.890 ;
        RECT  3.435 1.555 3.665 1.895 ;
        RECT  0.115 1.130 0.345 2.735 ;
        RECT  0.180 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.410 4.180 ;
        RECT  0.180 3.270 0.520 4.180 ;
        RECT  1.425 0.630 1.985 0.950 ;
        RECT  1.755 0.630 1.985 1.355 ;
        RECT  2.825 1.090 4.125 1.320 ;
        RECT  3.485 1.090 4.125 1.325 ;
        RECT  3.895 1.090 4.125 1.580 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  3.895 1.345 5.685 1.580 ;
        RECT  5.345 1.345 5.685 1.650 ;
        RECT  3.895 1.810 5.165 2.040 ;
        RECT  4.995 1.880 5.960 2.220 ;
        RECT  3.895 1.810 4.215 3.425 ;
        RECT  6.315 1.230 6.915 1.540 ;
        RECT  4.445 2.325 4.755 3.155 ;
        RECT  6.315 1.230 6.545 3.155 ;
        RECT  4.445 2.870 6.545 3.155 ;
        RECT  4.445 2.925 7.095 3.155 ;
        RECT  6.755 2.925 7.095 3.385 ;
        RECT  2.255 0.630 4.585 0.860 ;
        RECT  4.355 0.630 4.585 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.740 0.770 7.660 1.000 ;
        RECT  4.355 0.885 5.970 1.115 ;
        RECT  7.375 0.770 7.660 1.600 ;
        RECT  2.120 3.420 2.405 3.760 ;
        RECT  4.445 3.385 6.330 3.615 ;
        RECT  2.120 3.530 3.575 3.760 ;
        RECT  7.520 3.535 7.860 3.845 ;
        RECT  6.100 3.615 7.860 3.845 ;
        RECT  4.445 3.385 4.675 3.885 ;
        RECT  3.360 3.655 4.675 3.885 ;
        RECT  6.775 1.800 7.065 2.695 ;
        RECT  6.775 2.465 7.555 2.695 ;
        RECT  9.795 1.240 10.025 3.230 ;
        RECT  9.565 2.625 10.025 3.230 ;
        RECT  7.325 2.465 7.555 3.305 ;
        RECT  9.565 2.890 11.375 3.230 ;
        RECT  7.325 3.075 9.795 3.305 ;
        RECT  8.020 0.630 8.360 0.970 ;
        RECT  9.335 0.780 10.485 1.010 ;
        RECT  8.130 0.630 8.360 1.430 ;
        RECT  9.335 0.780 9.565 1.430 ;
        RECT  8.130 1.200 9.565 1.430 ;
        RECT  7.525 1.830 8.075 2.145 ;
        RECT  9.055 1.200 9.440 2.205 ;
        RECT  10.255 0.780 10.485 2.450 ;
        RECT  10.255 2.220 11.095 2.450 ;
        RECT  10.755 2.330 11.840 2.560 ;
        RECT  7.840 1.830 8.075 2.845 ;
        RECT  9.055 1.200 9.285 2.845 ;
        RECT  7.840 2.590 9.285 2.845 ;
        RECT  11.610 2.330 11.840 3.435 ;
        RECT  11.610 3.110 12.050 3.435 ;
        RECT  10.715 0.630 13.040 0.860 ;
        RECT  10.715 0.630 11.000 1.005 ;
        RECT  12.700 0.630 13.040 1.150 ;
        RECT  11.470 1.090 12.300 1.400 ;
        RECT  12.070 1.090 12.300 2.810 ;
        RECT  12.280 2.580 12.515 3.145 ;
        RECT  13.760 2.730 14.045 3.090 ;
        RECT  12.280 2.860 14.045 3.090 ;
        RECT  12.280 2.860 13.580 3.145 ;
        RECT  12.280 2.580 12.510 3.970 ;
        RECT  11.320 3.665 12.510 3.970 ;
        RECT  12.530 1.380 12.815 1.880 ;
        RECT  12.530 1.540 14.505 1.880 ;
        RECT  14.275 1.540 14.505 3.550 ;
        RECT  13.820 3.320 14.505 3.550 ;
        RECT  13.820 3.320 14.050 4.160 ;
        RECT  13.710 3.820 14.050 4.160 ;
        RECT  1.255 1.585 2.30 1.815 ;
        RECT  4.445 2.870 5.20 3.155 ;
        RECT  4.445 2.925 6.50 3.155 ;
        RECT  2.255 0.630 3.00 0.860 ;
        RECT  7.325 3.075 8.40 3.305 ;
        RECT  10.715 0.630 12.60 0.860 ;
    END
END SDFFRQX1

MACRO SDFFRQX0
    CLASS CORE ;
    FOREIGN SDFFRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.550  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.300 3.010 14.995 3.350 ;
        RECT  14.570 2.860 14.995 3.350 ;
        RECT  14.570 0.630 14.800 3.350 ;
        RECT  14.200 0.630 14.800 0.970 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.225 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.245 3.320 ;
        RECT  2.190 2.860 3.245 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.302  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.610 2.245 13.105 2.895 ;
        END
    END RN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.960 2.360 8.665 2.700 ;
        RECT  8.305 2.240 8.665 2.700 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.300 3.810 14.640 5.280 ;
        RECT  12.285 3.910 12.620 5.280 ;
        RECT  9.510 3.630 9.850 5.280 ;
        RECT  8.310 3.910 8.650 5.280 ;
        RECT  4.830 3.865 5.170 5.280 ;
        RECT  3.200 4.170 3.540 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.400 -0.400 13.740 0.950 ;
        RECT  8.615 -0.400 8.900 1.540 ;
        RECT  4.485 -0.400 4.825 0.655 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.270 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  0.750 0.630 1.675 0.950 ;
        RECT  1.445 0.630 1.675 1.355 ;
        RECT  1.445 1.125 3.730 1.355 ;
        RECT  3.185 1.090 3.730 1.355 ;
        RECT  3.500 1.345 5.425 1.575 ;
        RECT  3.505 1.805 5.520 2.090 ;
        RECT  5.235 1.805 5.520 2.180 ;
        RECT  3.505 1.805 3.735 3.480 ;
        RECT  3.505 3.140 4.140 3.480 ;
        RECT  5.750 1.230 6.655 1.540 ;
        RECT  3.965 2.325 4.950 2.665 ;
        RECT  4.605 2.325 4.950 3.175 ;
        RECT  4.605 2.945 5.980 3.175 ;
        RECT  5.750 1.230 5.980 3.175 ;
        RECT  5.805 3.025 6.500 3.230 ;
        RECT  5.830 3.025 6.500 3.255 ;
        RECT  6.270 3.025 6.500 3.790 ;
        RECT  6.270 3.450 6.610 3.790 ;
        RECT  4.370 3.405 5.625 3.635 ;
        RECT  4.370 3.405 4.600 3.940 ;
        RECT  1.995 3.710 4.600 3.940 ;
        RECT  5.420 3.430 5.650 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  7.030 3.910 7.370 4.250 ;
        RECT  5.420 4.020 7.370 4.250 ;
        RECT  1.980 0.630 4.190 0.860 ;
        RECT  3.960 0.630 4.190 1.115 ;
        RECT  1.980 0.630 2.320 0.895 ;
        RECT  5.290 0.770 7.455 1.000 ;
        RECT  3.960 0.885 5.520 1.115 ;
        RECT  7.115 0.770 7.455 1.570 ;
        RECT  6.210 2.510 7.075 2.795 ;
        RECT  9.590 1.230 9.820 3.330 ;
        RECT  8.080 2.990 10.800 3.330 ;
        RECT  10.455 2.990 10.800 3.395 ;
        RECT  6.845 2.510 7.075 3.680 ;
        RECT  8.080 2.990 8.310 3.680 ;
        RECT  6.845 3.450 8.310 3.680 ;
        RECT  9.130 0.770 10.280 1.000 ;
        RECT  7.815 1.230 8.155 2.010 ;
        RECT  7.815 1.780 9.360 2.010 ;
        RECT  6.495 1.800 9.360 2.010 ;
        RECT  9.130 0.770 9.360 2.010 ;
        RECT  6.210 1.840 8.045 2.110 ;
        RECT  6.210 1.840 7.730 2.180 ;
        RECT  10.050 0.770 10.280 2.425 ;
        RECT  10.050 2.195 10.800 2.425 ;
        RECT  10.460 2.305 11.595 2.535 ;
        RECT  8.895 1.780 9.235 2.650 ;
        RECT  7.500 1.800 7.730 3.220 ;
        RECT  7.500 2.925 7.825 3.220 ;
        RECT  7.500 2.930 7.850 3.220 ;
        RECT  11.255 2.305 11.595 3.440 ;
        RECT  10.510 0.635 12.860 0.865 ;
        RECT  12.520 0.635 12.860 0.970 ;
        RECT  10.510 0.635 10.850 0.975 ;
        RECT  11.485 1.175 12.055 1.515 ;
        RECT  12.805 3.125 13.610 3.465 ;
        RECT  11.825 3.235 13.610 3.465 ;
        RECT  10.805 3.640 11.140 3.970 ;
        RECT  10.805 3.655 11.145 3.970 ;
        RECT  11.825 1.175 12.055 3.970 ;
        RECT  10.805 3.685 12.055 3.970 ;
        RECT  13.840 1.410 14.340 1.750 ;
        RECT  12.450 1.695 14.070 2.015 ;
        RECT  13.840 1.410 14.070 4.175 ;
        RECT  13.195 3.835 14.070 4.175 ;
        RECT  0.980 1.585 2.50 1.960 ;
        RECT  1.445 1.125 2.10 1.355 ;
        RECT  3.505 1.805 4.40 2.090 ;
        RECT  1.995 3.710 3.60 3.940 ;
        RECT  1.980 0.630 3.40 0.860 ;
        RECT  5.290 0.770 6.80 1.000 ;
        RECT  8.080 2.990 9.40 3.330 ;
        RECT  6.495 1.800 8.40 2.010 ;
        RECT  10.510 0.635 11.30 0.865 ;
    END
END SDFFRQX0

MACRO SDFFQX4
    CLASS CORE ;
    FOREIGN SDFFQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 1.240 16.830 4.130 ;
        RECT  15.170 2.250 16.830 2.630 ;
        RECT  15.170 0.790 15.510 2.630 ;
        RECT  15.050 2.890 15.400 4.130 ;
        RECT  15.170 0.790 15.400 4.130 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.820 3.655 3.240 ;
        RECT  2.205 2.820 3.655 3.105 ;
        RECT  2.205 2.685 2.435 3.105 ;
        RECT  2.185 2.045 2.415 2.780 ;
        RECT  0.575 2.045 2.415 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.045 3.085 2.590 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.560 2.875 1.975 3.215 ;
        RECT  1.385 3.470 1.790 3.850 ;
        RECT  1.560 2.875 1.790 3.850 ;
        END
    END SD
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.135 1.640 8.695 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.930 -0.400 16.270 0.720 ;
        RECT  14.410 -0.400 14.750 0.710 ;
        RECT  13.005 -0.400 13.345 1.450 ;
        RECT  10.420 -0.400 10.760 1.370 ;
        RECT  8.415 -0.400 8.700 0.950 ;
        RECT  3.485 -0.400 4.935 0.710 ;
        RECT  1.425 -0.400 1.765 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 2.890 16.110 5.280 ;
        RECT  14.290 4.160 14.630 5.280 ;
        RECT  12.960 3.530 13.300 5.280 ;
        RECT  10.940 3.965 11.280 5.280 ;
        RECT  8.545 2.910 8.830 5.280 ;
        RECT  4.475 3.965 4.815 5.280 ;
        RECT  3.160 4.170 3.500 5.280 ;
        RECT  0.940 4.055 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.375 1.470 ;
        RECT  1.145 1.240 1.375 1.815 ;
        RECT  1.145 1.585 3.655 1.815 ;
        RECT  3.315 1.585 3.655 1.960 ;
        RECT  0.115 1.240 0.345 2.815 ;
        RECT  0.990 2.505 1.330 2.815 ;
        RECT  0.115 2.585 1.330 2.815 ;
        RECT  0.180 2.585 0.520 4.180 ;
        RECT  3.895 1.400 5.335 1.740 ;
        RECT  3.895 1.400 4.125 3.275 ;
        RECT  3.895 2.935 4.315 3.275 ;
        RECT  6.070 1.190 6.395 1.530 ;
        RECT  5.620 1.300 6.395 1.530 ;
        RECT  4.355 2.105 4.860 2.445 ;
        RECT  5.620 1.300 5.850 3.275 ;
        RECT  4.630 2.105 4.860 3.275 ;
        RECT  5.620 2.935 6.045 3.275 ;
        RECT  4.630 3.045 6.045 3.275 ;
        RECT  6.425 2.980 6.765 3.735 ;
        RECT  2.020 3.505 6.765 3.735 ;
        RECT  2.020 3.505 2.310 3.940 ;
        RECT  2.255 0.630 2.595 1.170 ;
        RECT  5.165 0.730 6.855 0.960 ;
        RECT  2.255 0.940 5.395 1.170 ;
        RECT  6.625 0.730 6.855 1.660 ;
        RECT  6.625 1.320 7.210 1.660 ;
        RECT  8.930 0.670 10.190 0.900 ;
        RECT  7.085 0.735 7.955 1.090 ;
        RECT  7.595 0.735 7.955 1.410 ;
        RECT  7.595 1.180 9.160 1.410 ;
        RECT  8.930 0.670 9.160 2.100 ;
        RECT  9.960 0.670 10.190 2.070 ;
        RECT  11.330 1.730 11.670 2.070 ;
        RECT  9.960 1.840 11.670 2.070 ;
        RECT  8.930 1.760 9.270 2.100 ;
        RECT  7.595 0.735 7.855 2.940 ;
        RECT  9.390 1.130 9.730 1.470 ;
        RECT  6.080 1.840 6.390 2.195 ;
        RECT  6.080 1.965 7.225 2.195 ;
        RECT  9.500 1.130 9.730 2.680 ;
        RECT  9.500 2.340 10.310 2.680 ;
        RECT  12.000 1.540 12.285 2.680 ;
        RECT  8.085 2.450 12.285 2.680 ;
        RECT  9.210 2.450 9.550 2.860 ;
        RECT  6.995 1.965 7.225 3.400 ;
        RECT  8.085 2.450 8.315 3.400 ;
        RECT  6.995 3.170 8.315 3.400 ;
        RECT  9.210 2.450 9.440 3.855 ;
        RECT  10.410 3.505 11.750 3.735 ;
        RECT  9.210 3.625 10.640 3.855 ;
        RECT  11.520 3.650 12.030 3.990 ;
        RECT  11.570 0.970 11.910 1.310 ;
        RECT  11.570 1.080 12.745 1.310 ;
        RECT  13.350 2.355 13.690 2.700 ;
        RECT  12.515 2.470 13.690 2.700 ;
        RECT  12.515 1.080 12.745 3.220 ;
        RECT  9.750 2.990 12.745 3.220 ;
        RECT  11.930 2.990 12.270 3.330 ;
        RECT  9.750 2.990 10.090 3.395 ;
        RECT  13.830 1.070 14.170 1.910 ;
        RECT  12.975 1.680 14.170 1.910 ;
        RECT  12.975 1.680 13.260 2.030 ;
        RECT  13.940 1.070 14.170 3.160 ;
        RECT  13.730 2.930 14.070 3.760 ;
        RECT  1.145 1.585 2.20 1.815 ;
        RECT  2.020 3.505 5.80 3.735 ;
        RECT  2.255 0.940 4.80 1.170 ;
        RECT  8.085 2.450 11.80 2.680 ;
        RECT  9.750 2.990 11.30 3.220 ;
    END
END SDFFQX4

MACRO SDFFQX2
    CLASS CORE ;
    FOREIGN SDFFQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.350 1.250 13.735 3.770 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.675 2.415 3.260 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.550 3.470 1.890 4.250 ;
        RECT  0.755 3.470 1.890 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.680 3.250 3.020 ;
        RECT  2.645 2.215 3.025 3.020 ;
        RECT  1.660 2.215 3.025 2.445 ;
        RECT  1.660 1.970 1.890 2.445 ;
        RECT  0.660 1.970 1.890 2.200 ;
        RECT  0.660 1.720 1.005 2.200 ;
        END
    END SE
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.515 2.250 8.065 2.630 ;
        RECT  7.515 2.020 7.800 2.630 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.910 -0.400 14.250 0.720 ;
        RECT  12.790 -0.400 13.130 0.720 ;
        RECT  11.385 -0.400 11.730 0.970 ;
        RECT  9.680 -0.400 10.020 0.790 ;
        RECT  7.560 -0.400 7.845 1.330 ;
        RECT  4.100 -0.400 4.440 0.710 ;
        RECT  2.800 -0.400 3.140 0.710 ;
        RECT  0.940 -0.400 1.280 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.910 4.170 14.250 5.280 ;
        RECT  12.795 4.170 13.135 5.280 ;
        RECT  11.185 3.960 11.525 5.280 ;
        RECT  9.005 3.660 9.345 5.280 ;
        RECT  7.705 3.530 8.045 5.280 ;
        RECT  4.415 4.100 4.755 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.080 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.035 0.520 1.420 ;
        RECT  0.180 1.190 1.540 1.420 ;
        RECT  1.310 1.190 1.540 1.740 ;
        RECT  1.310 1.510 3.060 1.740 ;
        RECT  2.720 1.510 3.060 1.985 ;
        RECT  0.180 1.035 0.410 4.110 ;
        RECT  0.180 2.430 1.360 2.660 ;
        RECT  1.020 2.430 1.360 2.770 ;
        RECT  0.180 2.430 0.520 4.110 ;
        RECT  3.480 1.400 3.840 2.015 ;
        RECT  3.480 1.785 5.160 2.015 ;
        RECT  4.890 1.785 5.160 2.485 ;
        RECT  3.480 1.400 3.710 3.240 ;
        RECT  3.480 2.900 4.200 3.240 ;
        RECT  5.330 1.205 5.670 1.545 ;
        RECT  3.940 2.245 4.660 2.585 ;
        RECT  4.430 2.245 4.660 2.945 ;
        RECT  4.430 2.715 5.620 2.945 ;
        RECT  5.390 1.205 5.620 3.385 ;
        RECT  5.390 3.045 5.985 3.385 ;
        RECT  1.770 0.630 2.110 1.170 ;
        RECT  4.690 0.745 6.470 0.975 ;
        RECT  1.770 0.940 4.920 1.170 ;
        RECT  6.130 0.745 6.470 1.595 ;
        RECT  6.405 3.530 6.745 3.870 ;
        RECT  2.120 3.640 6.745 3.870 ;
        RECT  2.120 3.640 2.410 4.020 ;
        RECT  8.075 0.630 9.450 0.860 ;
        RECT  6.785 0.630 7.125 0.965 ;
        RECT  9.220 0.630 9.450 1.920 ;
        RECT  6.895 1.560 8.305 1.790 ;
        RECT  8.075 0.630 8.305 1.890 ;
        RECT  9.220 1.690 10.550 1.920 ;
        RECT  10.210 1.690 10.550 2.030 ;
        RECT  8.295 1.660 8.530 2.120 ;
        RECT  6.895 0.630 7.125 2.165 ;
        RECT  6.520 1.825 7.285 2.165 ;
        RECT  6.945 1.560 7.285 2.825 ;
        RECT  8.535 1.090 8.990 1.430 ;
        RECT  5.850 1.900 6.190 2.625 ;
        RECT  5.850 2.395 6.445 2.625 ;
        RECT  9.675 2.360 11.060 2.700 ;
        RECT  8.760 2.470 11.060 2.700 ;
        RECT  6.215 2.395 6.445 3.300 ;
        RECT  8.465 2.960 8.990 3.300 ;
        RECT  8.760 1.090 8.990 3.300 ;
        RECT  6.215 3.055 8.990 3.300 ;
        RECT  10.560 0.630 10.900 0.970 ;
        RECT  10.670 0.630 10.900 1.460 ;
        RECT  10.670 1.230 11.520 1.460 ;
        RECT  11.290 1.230 11.520 3.160 ;
        RECT  12.370 2.340 12.655 3.160 ;
        RECT  10.155 2.930 12.655 3.160 ;
        RECT  10.155 2.930 10.495 3.825 ;
        RECT  12.090 0.680 12.430 2.105 ;
        RECT  11.750 1.875 13.115 2.105 ;
        RECT  11.750 1.875 12.040 2.650 ;
        RECT  12.885 1.875 13.115 3.730 ;
        RECT  12.030 3.390 13.115 3.730 ;
        RECT  1.770 0.940 3.70 1.170 ;
        RECT  2.120 3.640 5.30 3.870 ;
        RECT  8.760 2.470 10.70 2.700 ;
        RECT  6.215 3.055 7.10 3.300 ;
        RECT  10.155 2.930 11.30 3.160 ;
    END
END SDFFQX2

MACRO SDFFQX1
    CLASS CORE ;
    FOREIGN SDFFQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.420 2.250 14.375 2.630 ;
        RECT  13.160 3.780 13.650 4.120 ;
        RECT  13.420 0.700 13.650 4.120 ;
        RECT  13.160 0.700 13.650 1.040 ;
        END
    END Q
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 3.990 2.030 4.250 ;
        RECT  1.610 3.980 2.000 4.250 ;
        RECT  1.610 3.470 1.840 4.250 ;
        RECT  1.410 3.470 1.840 3.815 ;
        RECT  1.385 3.470 1.840 3.800 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.880 2.800 3.655 3.240 ;
        RECT  2.880 2.045 3.110 3.240 ;
        RECT  0.575 2.045 3.110 2.275 ;
        RECT  0.575 1.700 0.915 2.275 ;
        END
    END SE
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.580 2.650 3.190 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.640 8.225 2.085 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.880 3.330 14.220 5.280 ;
        RECT  12.365 4.040 12.705 5.280 ;
        RECT  9.480 3.500 9.820 5.280 ;
        RECT  8.180 3.620 8.520 5.280 ;
        RECT  4.905 3.845 5.230 5.280 ;
        RECT  3.260 4.170 3.600 5.280 ;
        RECT  0.940 4.005 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.880 -0.400 14.220 1.040 ;
        RECT  12.000 -0.400 12.340 1.050 ;
        RECT  10.145 -0.400 10.485 1.030 ;
        RECT  8.085 -0.400 8.425 0.950 ;
        RECT  4.725 -0.400 5.065 0.655 ;
        RECT  3.485 1.090 3.825 1.325 ;
        RECT  2.825 1.090 3.825 1.320 ;
        RECT  1.755 1.125 3.055 1.355 ;
        RECT  1.755 -0.400 1.985 1.355 ;
        RECT  1.425 -0.400 1.985 0.950 ;
        RECT  0.560 -0.400 0.900 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.560 1.130 0.900 1.470 ;
        RECT  0.115 1.240 1.485 1.470 ;
        RECT  1.255 1.240 1.485 1.815 ;
        RECT  1.255 1.585 3.630 1.815 ;
        RECT  3.290 1.555 3.630 1.895 ;
        RECT  0.115 1.240 0.345 2.790 ;
        RECT  0.115 2.505 1.360 2.790 ;
        RECT  0.180 2.505 0.520 4.180 ;
        RECT  3.900 1.755 4.240 2.110 ;
        RECT  3.900 1.880 5.275 2.110 ;
        RECT  4.935 1.880 5.275 2.220 ;
        RECT  3.900 1.755 4.215 3.425 ;
        RECT  5.885 1.200 6.225 1.540 ;
        RECT  4.445 2.565 4.775 3.155 ;
        RECT  5.680 1.310 5.920 3.155 ;
        RECT  4.445 2.925 6.460 3.155 ;
        RECT  6.120 2.925 6.460 3.460 ;
        RECT  2.255 0.630 4.495 0.860 ;
        RECT  4.265 0.630 4.495 1.115 ;
        RECT  2.255 0.630 2.595 0.895 ;
        RECT  5.295 0.740 6.995 0.970 ;
        RECT  4.265 0.885 5.525 1.115 ;
        RECT  6.685 0.740 6.995 1.685 ;
        RECT  2.070 3.420 2.410 3.760 ;
        RECT  4.445 3.385 5.710 3.615 ;
        RECT  5.480 3.385 5.710 3.930 ;
        RECT  2.070 3.530 3.580 3.760 ;
        RECT  4.445 3.385 4.675 3.885 ;
        RECT  3.365 3.655 4.675 3.885 ;
        RECT  6.880 3.620 7.220 3.930 ;
        RECT  5.480 3.700 7.220 3.930 ;
        RECT  9.115 1.095 9.455 1.460 ;
        RECT  6.165 2.165 6.505 2.675 ;
        RECT  6.165 2.445 6.995 2.675 ;
        RECT  9.115 1.095 9.345 3.230 ;
        RECT  8.940 2.710 9.345 3.230 ;
        RECT  6.765 2.445 6.995 3.390 ;
        RECT  8.940 2.890 10.730 3.230 ;
        RECT  6.765 3.160 9.170 3.390 ;
        RECT  8.655 0.630 9.915 0.860 ;
        RECT  7.225 0.645 7.625 1.410 ;
        RECT  8.655 0.630 8.885 1.410 ;
        RECT  7.225 1.180 8.885 1.410 ;
        RECT  8.485 1.180 8.820 1.980 ;
        RECT  6.965 1.915 7.455 2.205 ;
        RECT  9.685 0.630 9.915 2.450 ;
        RECT  9.685 2.220 10.465 2.450 ;
        RECT  10.125 2.330 11.210 2.560 ;
        RECT  7.225 0.645 7.455 2.930 ;
        RECT  7.225 2.690 7.760 2.930 ;
        RECT  10.980 2.330 11.210 3.320 ;
        RECT  10.980 2.980 11.405 3.320 ;
        RECT  10.995 0.705 11.670 1.070 ;
        RECT  11.440 2.430 11.885 2.660 ;
        RECT  11.440 0.705 11.670 2.660 ;
        RECT  11.650 2.660 12.520 3.000 ;
        RECT  10.630 3.545 10.930 3.840 ;
        RECT  10.740 3.550 10.970 4.215 ;
        RECT  11.650 2.430 11.880 4.215 ;
        RECT  10.740 3.985 11.880 4.215 ;
        RECT  11.900 1.615 13.140 1.955 ;
        RECT  11.900 1.615 12.185 2.135 ;
        RECT  12.910 1.615 13.140 3.470 ;
        RECT  12.460 3.240 13.140 3.470 ;
        RECT  12.460 3.240 12.800 3.580 ;
        RECT  1.255 1.585 2.20 1.815 ;
        RECT  4.445 2.925 5.80 3.155 ;
        RECT  2.255 0.630 3.60 0.860 ;
        RECT  6.765 3.160 8.60 3.390 ;
    END
END SDFFQX1

MACRO SDFFQX0
    CLASS CORE ;
    FOREIGN SDFFQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 1.640 13.105 2.020 ;
        RECT  12.620 3.430 12.960 3.770 ;
        RECT  12.725 1.640 12.960 3.770 ;
        RECT  12.725 0.630 12.955 3.770 ;
        RECT  12.045 0.630 12.955 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.190 3.215 2.630 ;
        END
    END D
    PIN SD
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 3.175 1.975 3.480 ;
        RECT  1.535 3.140 1.960 3.480 ;
        RECT  1.385 3.520 1.765 3.850 ;
        RECT  1.535 3.140 1.765 3.850 ;
        RECT  1.415 3.505 1.765 3.850 ;
        END
    END SD
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.239  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.905 2.860 3.215 3.320 ;
        RECT  2.190 2.860 3.215 3.090 ;
        RECT  2.185 2.250 2.415 3.020 ;
        RECT  2.015 2.250 2.415 2.640 ;
        RECT  0.705 2.250 2.415 2.550 ;
        END
    END SE
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.045 2.200 7.515 2.695 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  12.020 4.165 12.360 5.280 ;
        RECT  10.755 3.910 11.040 5.280 ;
        RECT  7.650 3.630 8.460 5.280 ;
        RECT  3.200 4.170 4.495 5.280 ;
        RECT  0.445 4.060 0.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  9.270 -0.400 9.555 0.710 ;
        RECT  9.250 -0.400 9.555 0.675 ;
        RECT  7.375 -0.400 7.660 0.970 ;
        RECT  3.970 -0.400 4.310 0.895 ;
        RECT  3.010 -0.400 3.350 0.710 ;
        RECT  0.750 -0.400 1.090 0.950 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.980 1.585 3.215 1.960 ;
        RECT  0.245 1.790 1.320 2.020 ;
        RECT  0.245 1.790 0.475 3.380 ;
        RECT  0.245 2.890 1.305 3.175 ;
        RECT  0.245 2.890 1.290 3.220 ;
        RECT  0.245 2.890 0.785 3.380 ;
        RECT  3.445 1.805 4.770 2.035 ;
        RECT  3.445 1.805 3.875 2.095 ;
        RECT  3.445 1.805 3.835 2.105 ;
        RECT  4.485 1.805 4.770 2.205 ;
        RECT  3.445 1.805 3.675 3.425 ;
        RECT  3.445 3.085 4.195 3.425 ;
        RECT  5.000 1.230 5.800 1.540 ;
        RECT  3.905 2.325 4.190 2.665 ;
        RECT  3.905 2.435 5.230 2.665 ;
        RECT  5.000 1.230 5.230 3.480 ;
        RECT  4.995 2.435 5.230 3.480 ;
        RECT  4.995 3.250 5.725 3.480 ;
        RECT  5.385 3.250 5.725 3.790 ;
        RECT  1.995 3.710 5.050 3.940 ;
        RECT  4.820 3.710 5.050 4.250 ;
        RECT  1.995 3.710 2.295 4.180 ;
        RECT  6.145 3.925 6.485 4.250 ;
        RECT  4.820 4.020 6.485 4.250 ;
        RECT  4.540 0.640 6.500 0.920 ;
        RECT  6.160 0.640 6.500 0.970 ;
        RECT  1.980 1.015 2.320 1.355 ;
        RECT  4.540 0.640 4.770 1.355 ;
        RECT  1.980 1.125 4.770 1.355 ;
        RECT  5.460 2.440 5.800 2.780 ;
        RECT  5.460 2.530 6.190 2.780 ;
        RECT  8.350 2.600 9.410 2.940 ;
        RECT  7.995 2.905 8.580 3.245 ;
        RECT  8.350 1.230 8.580 3.245 ;
        RECT  7.165 3.015 8.580 3.245 ;
        RECT  5.960 2.530 6.190 3.695 ;
        RECT  7.165 3.015 7.395 3.695 ;
        RECT  5.960 3.465 7.395 3.695 ;
        RECT  7.890 0.770 9.040 1.000 ;
        RECT  7.890 0.770 8.120 1.480 ;
        RECT  6.585 1.250 8.120 1.480 ;
        RECT  6.585 1.250 7.205 1.590 ;
        RECT  8.810 0.770 9.040 2.160 ;
        RECT  5.460 1.770 6.815 2.110 ;
        RECT  7.745 1.250 7.975 2.470 ;
        RECT  8.810 1.930 9.560 2.160 ;
        RECT  9.220 2.040 10.065 2.270 ;
        RECT  7.745 2.130 8.085 2.470 ;
        RECT  6.585 1.250 6.815 3.230 ;
        RECT  6.585 2.895 6.930 3.230 ;
        RECT  6.585 2.900 6.935 3.230 ;
        RECT  9.725 2.040 10.065 3.400 ;
        RECT  10.125 1.110 10.525 1.450 ;
        RECT  11.390 2.370 11.730 2.710 ;
        RECT  10.295 2.480 11.730 2.710 ;
        RECT  10.295 1.110 10.525 3.970 ;
        RECT  9.350 3.630 10.525 3.970 ;
        RECT  12.045 1.350 12.385 1.900 ;
        RECT  11.085 1.700 12.190 2.040 ;
        RECT  11.960 1.700 12.190 3.565 ;
        RECT  11.220 3.225 12.190 3.565 ;
        RECT  0.980 1.585 2.90 1.960 ;
        RECT  1.995 3.710 4.80 3.940 ;
        RECT  1.980 1.125 3.20 1.355 ;
    END
END SDFFQX0

MACRO OR8X1
    CLASS CORE ;
    FOREIGN OR8X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 1.690 1.765 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.660 1.640 1.135 2.485 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.250 7.580 2.630 ;
        RECT  7.240 1.670 7.580 2.630 ;
        END
    END B
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.745 3.120 2.030 ;
        RECT  2.780 1.695 3.115 2.030 ;
        RECT  2.780 1.030 3.025 2.030 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.365 3.790 4.025 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.476  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.620 2.240 6.185 2.640 ;
        RECT  5.720 2.240 6.060 3.790 ;
        RECT  5.620 0.720 5.960 2.660 ;
        RECT  4.280 2.430 6.060 2.660 ;
        RECT  4.280 2.430 4.620 3.810 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.345 1.605 6.955 2.025 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.845 1.860 8.245 2.210 ;
        RECT  7.685 2.860 8.125 3.250 ;
        RECT  7.845 1.860 8.125 3.250 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.640 2.435 2.380 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.360 -0.400 7.900 0.710 ;
        RECT  2.630 -0.400 4.320 0.745 ;
        RECT  0.980 -0.400 1.320 0.815 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.440 2.910 6.780 5.280 ;
        RECT  5.000 2.960 5.340 5.280 ;
        RECT  2.310 2.730 2.655 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.200 1.125 2.120 1.410 ;
        RECT  0.200 1.125 0.430 3.300 ;
        RECT  0.200 2.960 1.030 3.300 ;
        RECT  0.485 2.960 0.825 4.015 ;
        RECT  3.255 1.170 3.855 1.510 ;
        RECT  3.540 1.170 3.855 3.070 ;
        RECT  3.540 1.750 4.600 2.090 ;
        RECT  3.540 1.750 3.880 3.070 ;
        RECT  8.290 0.630 8.705 1.360 ;
        RECT  6.960 1.070 8.705 1.360 ;
        RECT  8.475 0.630 8.705 3.235 ;
        RECT  8.355 2.895 8.585 4.250 ;
        RECT  7.210 3.950 8.585 4.250 ;
    END
END OR8X1

MACRO OR8X0
    CLASS CORE ;
    FOREIGN OR8X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 1.685 1.135 2.275 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.300 1.645 6.950 1.875 ;
        RECT  6.300 1.615 6.925 1.910 ;
        RECT  6.300 1.615 6.825 2.025 ;
        RECT  6.300 1.540 6.805 2.025 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.290 1.670 7.630 2.010 ;
        RECT  7.290 1.670 7.520 2.580 ;
        RECT  7.055 2.100 7.435 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.895 1.670 8.245 2.010 ;
        RECT  7.685 2.750 8.125 3.240 ;
        RECT  7.895 1.670 8.125 3.240 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.685 2.435 2.350 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 1.885 1.765 2.630 ;
        END
    END E
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.745 3.120 2.030 ;
        RECT  2.780 1.695 3.115 2.030 ;
        RECT  2.780 1.030 3.025 2.030 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.275 3.790 4.025 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.658  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.910 2.730 6.250 3.070 ;
        RECT  5.715 2.235 6.195 2.745 ;
        RECT  4.310 2.205 6.000 2.435 ;
        RECT  5.660 0.960 6.000 2.435 ;
        RECT  4.310 2.205 4.650 3.070 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.360 -0.400 7.900 0.710 ;
        RECT  2.630 -0.400 4.320 0.745 ;
        RECT  0.980 -0.400 1.320 0.995 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.780 3.380 7.120 5.280 ;
        RECT  5.110 2.775 5.450 5.280 ;
        RECT  2.380 2.730 2.725 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.780 1.170 2.120 1.455 ;
        RECT  0.180 1.225 2.120 1.455 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  0.180 1.170 0.410 3.435 ;
        RECT  0.180 3.150 1.025 3.435 ;
        RECT  0.570 3.150 1.025 3.490 ;
        RECT  0.570 3.150 0.910 4.015 ;
        RECT  3.255 1.170 3.895 1.510 ;
        RECT  3.610 1.170 3.895 2.980 ;
        RECT  3.610 1.690 4.600 1.975 ;
        RECT  3.610 1.690 3.950 2.980 ;
        RECT  6.960 1.070 8.705 1.355 ;
        RECT  8.260 0.630 8.705 1.390 ;
        RECT  6.980 1.070 8.705 1.390 ;
        RECT  8.355 2.730 8.705 3.070 ;
        RECT  8.475 0.630 8.705 4.000 ;
        RECT  7.365 3.660 8.705 4.000 ;
    END
END OR8X0

MACRO OR7X1
    CLASS CORE ;
    FOREIGN OR7X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.345 1.585 6.990 2.025 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.476  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.620 2.240 6.195 2.640 ;
        RECT  5.720 2.240 6.060 3.790 ;
        RECT  5.620 0.720 5.960 2.730 ;
        RECT  4.280 2.500 6.060 2.730 ;
        RECT  4.280 2.500 4.620 3.810 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.275 3.790 4.025 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.745 3.120 2.030 ;
        RECT  2.780 1.695 3.115 2.030 ;
        RECT  2.780 1.030 3.025 2.030 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END G
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.660 1.640 1.135 2.510 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.640 2.435 2.380 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.250 7.615 2.665 ;
        RECT  7.330 1.670 7.615 2.665 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 1.690 1.765 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.440 2.910 6.780 5.280 ;
        RECT  5.000 2.960 5.340 5.280 ;
        RECT  2.310 2.730 2.655 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.360 -0.400 7.900 0.710 ;
        RECT  2.630 -0.400 4.320 0.745 ;
        RECT  0.980 -0.400 1.320 0.815 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.200 1.125 2.120 1.410 ;
        RECT  0.200 1.125 0.430 3.300 ;
        RECT  0.200 2.960 1.030 3.300 ;
        RECT  0.485 2.960 0.825 4.015 ;
        RECT  3.255 1.170 3.895 1.510 ;
        RECT  3.580 1.170 3.895 2.980 ;
        RECT  3.580 1.750 4.600 2.090 ;
        RECT  3.580 1.750 3.920 2.980 ;
        RECT  6.960 1.070 8.075 1.355 ;
        RECT  7.845 1.070 8.075 3.235 ;
        RECT  7.670 2.910 7.900 4.150 ;
        RECT  7.210 3.810 7.900 4.150 ;
    END
END OR7X1

MACRO OR7X0
    CLASS CORE ;
    FOREIGN OR7X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.658  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.840 2.235 6.195 3.065 ;
        RECT  5.660 0.960 6.000 2.640 ;
        RECT  4.310 2.410 6.195 2.640 ;
        RECT  4.310 2.410 4.650 3.065 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.270 3.740 3.930 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.745 3.120 2.030 ;
        RECT  2.780 1.695 3.115 2.030 ;
        RECT  2.780 1.030 3.025 2.030 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.090 1.765 3.265 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.685 2.435 2.380 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.290 1.670 7.615 2.445 ;
        RECT  7.055 2.230 7.495 2.660 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.300 1.640 6.950 1.985 ;
        RECT  6.300 1.640 6.805 2.025 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 1.690 1.135 2.735 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.640 3.375 6.980 5.280 ;
        RECT  5.040 3.370 5.380 5.280 ;
        RECT  2.380 2.730 2.725 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.360 -0.400 7.900 0.710 ;
        RECT  2.630 -0.400 4.320 0.745 ;
        RECT  0.980 -0.400 1.320 0.995 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.780 1.170 2.120 1.455 ;
        RECT  0.180 1.225 2.120 1.455 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  0.240 1.170 0.470 3.430 ;
        RECT  0.240 3.145 1.025 3.430 ;
        RECT  0.570 3.145 1.025 3.485 ;
        RECT  0.570 3.145 0.910 4.010 ;
        RECT  3.255 1.170 3.895 1.510 ;
        RECT  3.610 1.170 3.895 2.980 ;
        RECT  3.610 1.690 4.600 2.030 ;
        RECT  3.610 1.690 3.950 2.980 ;
        RECT  6.960 1.070 8.075 1.390 ;
        RECT  7.845 1.070 8.075 3.065 ;
        RECT  7.720 2.725 7.950 3.995 ;
        RECT  7.365 3.655 7.950 3.995 ;
    END
END OR7X0

MACRO OR6X4
    CLASS CORE ;
    FOREIGN OR6X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.590 1.430 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.750 4.000 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 0.890 10.585 3.895 ;
        RECT  8.790 2.050 10.585 2.280 ;
        RECT  8.750 2.640 9.090 3.900 ;
        RECT  8.790 0.890 9.090 3.900 ;
        RECT  8.750 0.890 9.090 1.700 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.880 5.940 2.220 ;
        RECT  5.165 1.640 5.560 2.220 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.640 6.775 1.990 ;
        RECT  6.270 1.660 6.755 2.020 ;
        RECT  6.270 1.660 6.735 2.220 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 3.470 2.530 4.000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.335 2.250 1.880 2.700 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 2.640 9.810 5.280 ;
        RECT  7.990 2.640 8.330 5.280 ;
        RECT  5.360 3.065 5.700 5.280 ;
        RECT  3.860 3.225 4.200 5.280 ;
        RECT  1.370 3.900 1.710 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.700 ;
        RECT  8.030 -0.400 8.370 1.700 ;
        RECT  6.610 -0.400 6.950 0.840 ;
        RECT  5.190 -0.400 5.530 1.410 ;
        RECT  2.810 -0.400 3.150 0.710 ;
        RECT  1.580 -0.400 1.920 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.210 1.400 2.565 2.265 ;
        RECT  2.420 1.930 3.505 2.270 ;
        RECT  2.420 1.930 2.770 3.200 ;
        RECT  1.580 0.940 4.570 1.170 ;
        RECT  0.115 1.020 1.810 1.360 ;
        RECT  4.340 0.940 4.570 2.530 ;
        RECT  4.340 2.190 4.680 2.530 ;
        RECT  0.115 1.020 0.345 3.240 ;
        RECT  0.115 2.890 0.520 3.240 ;
        RECT  5.990 0.630 6.330 1.430 ;
        RECT  6.510 2.910 6.850 4.250 ;
        RECT  6.240 3.950 6.850 4.250 ;
        RECT  3.510 1.400 4.035 1.700 ;
        RECT  6.965 2.120 7.280 2.460 ;
        RECT  4.910 2.450 7.195 2.680 ;
        RECT  3.735 1.400 4.035 2.995 ;
        RECT  4.910 2.450 5.140 2.990 ;
        RECT  3.140 2.760 4.920 2.995 ;
        RECT  3.140 2.760 3.480 3.700 ;
        RECT  4.580 2.760 4.920 3.700 ;
        RECT  7.310 0.700 7.740 1.700 ;
        RECT  7.510 1.945 8.560 2.285 ;
        RECT  7.510 0.700 7.740 4.180 ;
        RECT  7.270 2.915 7.740 4.180 ;
        RECT  1.580 0.940 3.80 1.170 ;
        RECT  4.910 2.450 6.30 2.680 ;
    END
END OR6X4

MACRO OR6X2
    CLASS CORE ;
    FOREIGN OR6X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.570 0.585 2.100 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.650 1.640 8.070 2.225 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.695 2.120 3.350 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.120 2.465 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 1.760 8.735 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.035 3.010 7.375 3.880 ;
        RECT  5.210 3.010 7.375 3.305 ;
        RECT  5.555 3.010 5.895 3.880 ;
        RECT  5.215 1.525 5.895 1.870 ;
        RECT  5.555 1.000 5.895 1.870 ;
        RECT  4.115 3.080 5.895 3.310 ;
        RECT  5.210 2.900 5.545 3.310 ;
        RECT  5.215 1.525 5.545 3.310 ;
        RECT  4.115 3.080 4.455 3.880 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.275 2.120 1.765 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.780 3.320 8.120 5.280 ;
        RECT  6.275 3.540 6.615 5.280 ;
        RECT  4.835 3.540 5.175 5.280 ;
        RECT  3.355 3.320 3.700 5.280 ;
        RECT  0.175 2.640 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.655 -0.400 8.995 0.950 ;
        RECT  7.135 -0.400 7.475 1.445 ;
        RECT  3.725 -0.400 4.065 0.970 ;
        RECT  1.620 -0.400 2.440 1.430 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.150 1.240 1.890 ;
        RECT  0.815 1.660 4.315 1.890 ;
        RECT  3.975 1.660 4.315 2.390 ;
        RECT  0.815 1.660 1.045 3.090 ;
        RECT  0.815 2.860 1.670 3.090 ;
        RECT  1.330 2.860 1.670 3.960 ;
        RECT  2.965 1.090 3.305 1.430 ;
        RECT  2.965 1.200 4.985 1.430 ;
        RECT  4.645 1.200 4.985 2.850 ;
        RECT  3.580 2.620 4.985 2.850 ;
        RECT  3.580 2.620 3.810 3.090 ;
        RECT  2.100 2.860 3.810 3.090 ;
        RECT  2.100 2.860 2.440 3.960 ;
        RECT  7.895 1.060 8.235 1.410 ;
        RECT  7.895 1.180 9.270 1.410 ;
        RECT  5.795 2.440 6.135 2.780 ;
        RECT  5.795 2.550 8.010 2.780 ;
        RECT  7.780 2.550 8.010 3.090 ;
        RECT  7.780 2.860 9.270 3.090 ;
        RECT  9.015 1.180 9.270 3.960 ;
        RECT  8.930 2.855 9.270 3.960 ;
        RECT  0.815 1.660 3.70 1.890 ;
        RECT  2.965 1.200 3.30 1.430 ;
        RECT  5.795 2.550 7.70 2.780 ;
    END
END OR6X2

MACRO OR6X1
    CLASS CORE ;
    FOREIGN OR6X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 1.640 1.135 2.020 ;
        RECT  0.575 1.640 0.915 2.120 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.393  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.540 4.935 3.810 ;
        RECT  4.440 0.720 4.780 2.770 ;
        RECT  3.205 2.540 4.935 2.770 ;
        RECT  3.205 2.540 3.490 3.750 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.250 6.355 2.630 ;
        RECT  6.020 1.690 6.355 2.630 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.940 1.780 2.395 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.345 3.470 2.975 3.870 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.030 1.765 1.410 ;
        RECT  1.270 2.210 1.615 2.550 ;
        RECT  1.385 1.030 1.615 2.550 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.040 1.640 5.680 2.030 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.350 3.660 5.690 5.280 ;
        RECT  3.870 3.000 4.210 5.280 ;
        RECT  1.435 2.870 1.775 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.140 -0.400 6.680 0.710 ;
        RECT  1.620 -0.400 3.160 0.800 ;
        RECT  0.220 -0.400 0.560 0.770 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.820 1.070 1.155 1.410 ;
        RECT  0.115 1.180 1.155 1.410 ;
        RECT  0.115 1.180 0.345 4.250 ;
        RECT  0.115 2.870 0.600 3.210 ;
        RECT  0.115 2.870 0.505 4.250 ;
        RECT  2.220 1.210 2.950 1.550 ;
        RECT  2.720 1.995 3.440 2.310 ;
        RECT  2.720 1.210 2.950 3.070 ;
        RECT  2.610 2.730 2.950 3.070 ;
        RECT  5.740 1.070 6.815 1.410 ;
        RECT  6.410 2.860 6.815 3.200 ;
        RECT  6.585 1.070 6.815 4.250 ;
        RECT  5.920 3.910 6.815 4.250 ;
    END
END OR6X1

MACRO OR6X0
    CLASS CORE ;
    FOREIGN OR6X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.250 6.355 2.630 ;
        RECT  6.070 1.855 6.355 2.630 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.145 2.250 1.765 2.630 ;
        RECT  1.145 1.850 1.435 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.640 0.455 2.250 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.900 1.640 2.450 2.030 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.235 3.470 3.025 3.850 ;
        RECT  2.235 3.275 2.580 3.850 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.737  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.730 4.915 3.070 ;
        RECT  4.510 2.250 4.915 3.070 ;
        RECT  4.510 0.960 4.865 3.070 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.590 5.730 2.025 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.380 3.380 5.720 5.280 ;
        RECT  3.780 3.380 4.120 5.280 ;
        RECT  1.445 3.410 1.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.210 -0.400 6.750 0.710 ;
        RECT  1.580 -0.400 3.190 0.710 ;
        RECT  0.245 -0.400 0.585 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.685 1.170 1.025 1.510 ;
        RECT  0.685 1.170 0.915 3.075 ;
        RECT  0.180 2.730 0.915 3.075 ;
        RECT  0.180 2.730 0.520 4.015 ;
        RECT  2.180 1.070 2.975 1.410 ;
        RECT  2.715 1.070 2.975 1.975 ;
        RECT  2.715 1.690 3.470 1.975 ;
        RECT  2.715 1.070 2.945 2.980 ;
        RECT  2.475 2.640 2.945 2.980 ;
        RECT  5.810 1.070 6.815 1.370 ;
        RECT  6.585 1.070 6.815 4.000 ;
        RECT  6.425 2.895 6.815 4.000 ;
    END
END OR6X0

MACRO OR5X4
    CLASS CORE ;
    FOREIGN OR5X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.380 4.250 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.585 2.640 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 0.890 9.325 3.895 ;
        RECT  7.530 2.050 9.325 2.280 ;
        RECT  7.490 2.640 7.830 3.900 ;
        RECT  7.530 0.890 7.830 3.900 ;
        RECT  7.490 0.890 7.830 1.700 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.590 2.070 2.020 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.470 3.170 4.000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.970 2.250 2.515 2.695 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.210 2.640 8.550 5.280 ;
        RECT  6.730 2.640 7.070 5.280 ;
        RECT  4.490 3.225 4.830 5.280 ;
        RECT  1.860 2.975 2.200 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.210 -0.400 8.550 1.700 ;
        RECT  6.770 -0.400 7.110 1.700 ;
        RECT  4.095 -0.400 4.435 1.315 ;
        RECT  2.380 -0.400 2.720 0.710 ;
        RECT  0.990 -0.400 1.330 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.380 0.940 3.865 1.170 ;
        RECT  0.115 1.020 2.610 1.360 ;
        RECT  3.635 0.940 3.865 2.070 ;
        RECT  3.635 1.730 4.590 2.070 ;
        RECT  0.825 1.020 1.055 3.240 ;
        RECT  0.220 2.890 1.055 3.240 ;
        RECT  3.060 1.400 3.405 3.200 ;
        RECT  4.960 2.190 5.310 2.530 ;
        RECT  3.060 2.300 5.310 2.530 ;
        RECT  3.060 2.300 3.410 3.200 ;
        RECT  5.215 1.050 5.770 1.390 ;
        RECT  5.540 2.120 6.020 2.460 ;
        RECT  5.540 1.050 5.770 2.990 ;
        RECT  3.770 2.760 5.550 2.995 ;
        RECT  3.770 2.760 4.110 3.700 ;
        RECT  5.210 2.760 5.550 3.700 ;
        RECT  6.050 0.700 6.480 1.700 ;
        RECT  6.250 1.945 7.300 2.285 ;
        RECT  6.250 0.700 6.480 4.180 ;
        RECT  6.010 2.690 6.480 4.180 ;
        RECT  0.115 1.020 1.90 1.360 ;
        RECT  3.060 2.300 4.70 2.530 ;
    END
END OR5X4

MACRO OR5X2
    CLASS CORE ;
    FOREIGN OR5X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.615 2.345 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.315 2.860 1.765 3.240 ;
        RECT  1.315 2.120 1.715 3.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.120 1.085 2.685 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.845 1.800 6.345 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.501  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.375 3.035 4.715 3.960 ;
        RECT  2.935 3.035 4.715 3.330 ;
        RECT  3.275 2.860 3.870 3.330 ;
        RECT  3.530 1.170 3.870 3.330 ;
        RECT  2.935 3.035 3.275 3.960 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 2.120 2.385 2.685 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.095 3.320 5.435 5.280 ;
        RECT  3.655 3.560 3.995 5.280 ;
        RECT  2.175 2.915 2.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.285 -0.400 6.625 0.950 ;
        RECT  4.680 -0.400 5.020 1.455 ;
        RECT  2.380 -0.400 2.720 1.430 ;
        RECT  0.900 -0.400 1.240 1.430 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.130 0.520 1.890 ;
        RECT  1.620 1.180 1.960 1.890 ;
        RECT  0.115 1.660 2.955 1.890 ;
        RECT  2.615 1.660 2.955 2.220 ;
        RECT  0.115 1.130 0.345 4.180 ;
        RECT  0.115 2.915 0.520 4.180 ;
        RECT  5.525 1.060 5.865 1.410 ;
        RECT  5.525 1.180 6.805 1.410 ;
        RECT  4.135 2.465 4.475 2.805 ;
        RECT  4.135 2.575 5.615 2.805 ;
        RECT  5.385 2.575 5.615 3.090 ;
        RECT  5.385 2.860 6.805 3.090 ;
        RECT  6.575 1.180 6.805 3.960 ;
        RECT  6.370 2.860 6.805 3.960 ;
        RECT  0.115 1.660 1.80 1.890 ;
    END
END OR5X2

MACRO OR5X1
    CLASS CORE ;
    FOREIGN OR5X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.680 2.250 1.135 2.785 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.964  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 0.990 3.610 1.330 ;
        RECT  3.180 2.255 3.520 3.360 ;
        RECT  2.810 2.255 3.520 2.485 ;
        RECT  2.810 0.990 3.040 2.485 ;
        RECT  2.645 0.990 3.040 1.410 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.940 1.945 2.395 2.685 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.810 1.690 5.095 2.390 ;
        RECT  4.535 2.860 4.975 3.240 ;
        RECT  4.745 2.160 4.975 3.240 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.130 1.660 4.470 2.030 ;
        RECT  3.275 1.640 4.395 2.025 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 2.860 1.765 3.240 ;
        RECT  1.365 1.645 1.595 3.240 ;
        RECT  1.235 1.645 1.595 1.985 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.085 -0.400 5.445 0.710 ;
        RECT  0.925 -0.400 2.380 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.920 3.130 4.260 5.280 ;
        RECT  2.420 3.020 2.765 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.415 ;
        RECT  0.180 1.110 1.820 1.415 ;
        RECT  0.180 3.020 0.735 3.360 ;
        RECT  0.180 0.630 0.435 4.250 ;
        RECT  0.180 3.910 0.545 4.250 ;
        RECT  4.605 1.170 5.555 1.460 ;
        RECT  5.205 2.980 5.555 3.320 ;
        RECT  5.325 1.170 5.555 4.250 ;
        RECT  4.690 3.950 5.555 4.250 ;
    END
END OR5X1

MACRO OR5X0
    CLASS CORE ;
    FOREIGN OR5X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.640 1.730 1.135 2.630 ;
        RECT  0.685 1.720 1.135 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.690 4.470 2.030 ;
        RECT  3.275 1.640 3.655 2.030 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.810 1.690 5.095 2.390 ;
        RECT  4.535 2.860 4.975 3.240 ;
        RECT  4.745 2.185 4.975 3.240 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 1.720 2.425 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 2.860 1.765 3.240 ;
        RECT  1.365 1.720 1.650 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.619  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.320 2.300 3.660 3.360 ;
        RECT  2.815 0.630 3.550 0.930 ;
        RECT  2.815 2.300 3.660 2.530 ;
        RECT  2.815 0.630 3.045 2.530 ;
        RECT  2.645 1.030 3.045 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.120 3.670 4.460 5.280 ;
        RECT  2.400 3.020 2.745 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.950 -0.400 5.490 0.710 ;
        RECT  0.980 -0.400 2.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 1.920 1.455 ;
        RECT  1.580 1.170 1.920 1.460 ;
        RECT  0.180 1.170 0.515 1.505 ;
        RECT  0.180 1.170 0.410 3.325 ;
        RECT  0.180 3.020 0.925 3.325 ;
        RECT  0.470 3.020 0.925 3.360 ;
        RECT  0.470 3.020 0.810 3.940 ;
        RECT  4.550 1.170 5.555 1.460 ;
        RECT  5.205 3.020 5.555 3.360 ;
        RECT  5.325 1.170 5.555 4.250 ;
        RECT  4.690 3.950 5.555 4.250 ;
    END
END OR5X0

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.590 1.430 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.750 4.000 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 0.890 8.695 3.895 ;
        RECT  6.900 2.050 8.695 2.280 ;
        RECT  6.860 2.640 7.200 3.900 ;
        RECT  6.900 0.890 7.200 3.900 ;
        RECT  6.860 0.890 7.200 1.700 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 3.470 2.530 4.000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.335 2.250 1.880 2.700 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 2.640 7.920 5.280 ;
        RECT  6.100 2.640 6.440 5.280 ;
        RECT  3.860 3.225 4.200 5.280 ;
        RECT  1.370 3.900 1.710 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.700 ;
        RECT  6.140 -0.400 6.480 1.700 ;
        RECT  4.720 -0.400 5.060 1.705 ;
        RECT  2.810 -0.400 3.150 0.710 ;
        RECT  1.580 -0.400 1.920 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.210 1.400 2.565 2.265 ;
        RECT  2.420 1.930 3.505 2.270 ;
        RECT  2.420 1.930 2.770 3.200 ;
        RECT  1.580 0.940 4.445 1.170 ;
        RECT  0.115 1.020 1.810 1.360 ;
        RECT  4.215 0.940 4.445 2.530 ;
        RECT  4.215 2.190 4.680 2.530 ;
        RECT  0.115 1.020 0.345 3.240 ;
        RECT  0.115 2.890 0.520 3.240 ;
        RECT  3.510 1.400 3.985 1.700 ;
        RECT  5.050 2.120 5.390 2.460 ;
        RECT  4.910 2.450 5.305 2.680 ;
        RECT  3.735 1.400 3.985 2.995 ;
        RECT  4.910 2.450 5.140 2.990 ;
        RECT  3.140 2.760 4.920 2.995 ;
        RECT  3.140 2.760 3.480 3.700 ;
        RECT  4.580 2.760 4.920 3.700 ;
        RECT  5.420 0.700 5.850 1.700 ;
        RECT  5.620 1.945 6.670 2.285 ;
        RECT  5.620 0.700 5.850 4.180 ;
        RECT  5.380 2.915 5.850 4.180 ;
        RECT  1.580 0.940 3.30 1.170 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.640 4.940 2.230 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.315 2.120 1.755 2.685 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.120 1.085 2.685 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.170 1.880 5.660 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.526  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.665 3.035 4.005 3.960 ;
        RECT  2.225 3.035 4.005 3.330 ;
        RECT  2.645 2.860 3.235 3.330 ;
        RECT  2.895 1.170 3.235 3.330 ;
        RECT  2.225 3.035 2.565 3.960 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.410 3.320 4.750 5.280 ;
        RECT  2.945 3.560 3.285 5.280 ;
        RECT  1.435 2.915 1.780 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.600 -0.400 5.940 0.950 ;
        RECT  4.045 -0.400 4.385 1.455 ;
        RECT  1.660 -0.400 2.000 1.430 ;
        RECT  0.180 -0.400 0.520 1.430 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.180 1.240 1.890 ;
        RECT  0.115 1.660 2.325 1.890 ;
        RECT  1.985 1.660 2.325 2.220 ;
        RECT  0.115 1.660 0.345 3.960 ;
        RECT  0.115 2.915 0.520 3.960 ;
        RECT  4.840 1.060 5.220 1.410 ;
        RECT  4.840 1.180 6.120 1.410 ;
        RECT  3.465 2.465 3.805 2.805 ;
        RECT  3.465 2.575 4.640 2.805 ;
        RECT  4.410 2.575 4.640 3.090 ;
        RECT  4.410 2.860 6.120 3.090 ;
        RECT  5.890 1.180 6.120 3.960 ;
        RECT  5.740 2.855 6.120 3.960 ;
        RECT  0.115 1.660 1.20 1.890 ;
    END
END OR4X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.840 2.025 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.310 1.945 1.765 2.685 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.695 2.860 1.135 3.240 ;
        RECT  0.695 1.690 0.925 3.240 ;
        RECT  0.575 1.690 0.925 2.030 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.180 1.670 4.465 2.390 ;
        RECT  3.905 2.860 4.345 3.240 ;
        RECT  4.115 2.160 4.345 3.240 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.992  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 0.990 2.960 1.330 ;
        RECT  2.550 2.255 2.890 3.360 ;
        RECT  2.180 2.255 2.890 2.485 ;
        RECT  2.180 0.990 2.410 2.485 ;
        RECT  2.015 0.990 2.410 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.290 3.130 3.630 5.280 ;
        RECT  1.790 3.020 2.135 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.400 -0.400 4.860 0.710 ;
        RECT  0.180 -0.400 1.635 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.170 1.125 1.460 ;
        RECT  0.115 3.020 0.465 3.360 ;
        RECT  0.115 1.170 0.345 4.250 ;
        RECT  0.115 3.910 0.505 4.250 ;
        RECT  3.920 1.110 4.925 1.415 ;
        RECT  3.935 1.110 4.925 1.430 ;
        RECT  4.575 2.980 4.925 3.320 ;
        RECT  4.695 1.110 4.925 4.250 ;
        RECT  4.060 3.950 4.925 4.250 ;
    END
END OR4X1

MACRO OR4X0
    CLASS CORE ;
    FOREIGN OR4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.840 2.025 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.180 1.670 4.465 2.390 ;
        RECT  3.905 2.860 4.345 3.240 ;
        RECT  4.115 2.160 4.345 3.240 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.310 1.945 1.765 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.695 2.860 1.135 3.240 ;
        RECT  0.695 1.690 0.980 3.240 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.619  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.690 2.255 3.030 3.360 ;
        RECT  2.180 0.630 2.850 0.930 ;
        RECT  2.180 2.255 3.030 2.485 ;
        RECT  2.180 0.630 2.410 2.485 ;
        RECT  2.015 1.030 2.410 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.490 3.670 3.830 5.280 ;
        RECT  1.770 3.020 2.115 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.210 -0.400 4.750 0.710 ;
        RECT  0.180 -0.400 1.795 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 1.195 1.460 ;
        RECT  0.180 1.170 0.465 4.040 ;
        RECT  0.180 3.700 0.610 4.040 ;
        RECT  3.810 1.070 4.925 1.410 ;
        RECT  4.575 3.020 4.925 3.360 ;
        RECT  4.695 1.070 4.925 4.250 ;
        RECT  4.060 3.950 4.925 4.250 ;
    END
END OR4X0

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.135 1.640 6.805 2.220 ;
        RECT  2.975 1.640 6.805 1.890 ;
        RECT  2.975 1.640 3.315 2.460 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.460 2.120 5.805 2.460 ;
        RECT  3.955 2.860 5.690 3.090 ;
        RECT  5.460 2.120 5.690 3.090 ;
        RECT  3.955 2.120 4.285 3.090 ;
        RECT  3.935 2.120 4.285 2.595 ;
        RECT  3.645 2.120 4.285 2.460 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.120 4.995 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 1.350 1.960 3.895 ;
        RECT  0.125 1.930 1.960 2.330 ;
        RECT  0.125 0.700 0.520 3.895 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 0.710 ;
        RECT  5.215 -0.400 5.560 0.710 ;
        RECT  3.700 -0.400 4.040 0.950 ;
        RECT  2.180 -0.400 2.520 0.710 ;
        RECT  0.900 -0.400 1.240 1.700 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.380 2.640 6.720 5.280 ;
        RECT  2.540 3.150 2.880 5.280 ;
        RECT  0.900 2.635 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.940 1.050 3.280 1.410 ;
        RECT  2.190 1.160 3.280 1.410 ;
        RECT  4.460 1.050 4.800 1.410 ;
        RECT  5.780 1.120 6.120 1.410 ;
        RECT  2.190 1.180 6.120 1.410 ;
        RECT  2.190 1.160 2.530 2.920 ;
        RECT  2.190 2.690 3.725 2.920 ;
        RECT  3.495 2.690 3.725 3.550 ;
        RECT  3.495 3.320 4.895 3.550 ;
        RECT  4.555 3.320 4.895 4.180 ;
        RECT  2.190 1.180 5.80 1.410 ;
    END
END OR3X4

MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 2.290 2.355 2.630 ;
        RECT  1.905 2.080 2.345 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.275 2.860 1.765 3.240 ;
        RECT  1.275 2.120 1.615 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.585 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.295 1.660 3.640 2.020 ;
        RECT  3.295 1.640 3.605 2.020 ;
        RECT  3.295 1.210 3.525 2.965 ;
        RECT  2.975 2.640 3.360 3.560 ;
        RECT  3.035 1.210 3.525 1.550 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.755 2.640 4.095 5.280 ;
        RECT  2.225 2.860 2.565 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.755 -0.400 4.095 1.460 ;
        RECT  2.265 -0.400 2.605 1.240 ;
        RECT  0.740 -0.400 1.080 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.120 0.520 1.410 ;
        RECT  0.180 1.180 1.045 1.410 ;
        RECT  0.815 1.360 1.845 1.700 ;
        RECT  0.815 1.470 2.805 1.700 ;
        RECT  2.575 1.470 2.805 2.220 ;
        RECT  2.575 1.880 3.065 2.220 ;
        RECT  0.815 1.180 1.045 2.870 ;
        RECT  0.180 2.640 1.045 2.870 ;
        RECT  0.180 2.640 0.520 4.180 ;
    END
END OR3X2

MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.520 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.080 1.785 2.690 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.120 0.695 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.220 2.860 3.665 3.240 ;
        RECT  3.435 1.120 3.665 3.240 ;
        RECT  3.220 1.120 3.665 1.460 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.460 3.740 2.800 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.460 -0.400 2.800 1.065 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.240 0.520 1.580 ;
        RECT  1.660 1.240 2.000 1.580 ;
        RECT  0.180 1.350 2.990 1.580 ;
        RECT  2.760 1.350 2.990 2.220 ;
        RECT  2.760 1.880 3.190 2.220 ;
        RECT  0.925 1.350 1.155 3.155 ;
        RECT  0.180 2.925 1.155 3.155 ;
        RECT  0.180 2.925 0.520 3.265 ;
        RECT  0.180 1.350 1.60 1.580 ;
    END
END OR3X1

MACRO OR3X0
    CLASS CORE ;
    FOREIGN OR3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.540 1.920 2.125 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.155 2.630 ;
        RECT  0.870 1.690 1.155 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.540 0.505 2.225 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.558  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.495 2.860 3.035 3.380 ;
        RECT  2.805 0.630 3.035 3.380 ;
        RECT  2.630 0.630 3.035 0.970 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.640 3.690 1.980 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.930 -0.400 2.270 0.720 ;
        RECT  0.460 -0.400 0.800 1.265 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.330 1.025 2.380 1.310 ;
        RECT  2.150 1.025 2.380 2.545 ;
        RECT  2.150 2.205 2.575 2.545 ;
        RECT  2.035 2.340 2.265 3.380 ;
        RECT  0.180 3.040 2.265 3.380 ;
        RECT  0.180 3.040 1.40 3.380 ;
    END
END OR3X0

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.827  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.280 2.860 4.850 3.240 ;
        RECT  3.650 1.440 3.885 3.240 ;
        RECT  3.380 0.700 3.720 1.785 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.742  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.870 2.590 2.210 ;
        RECT  0.420 2.440 2.395 2.670 ;
        RECT  2.015 1.870 2.395 2.670 ;
        RECT  0.420 1.870 0.760 2.670 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.742  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.355 1.640 1.785 2.210 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.150 -0.400 4.490 1.685 ;
        RECT  2.620 -0.400 2.960 0.710 ;
        RECT  1.500 -0.400 1.840 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.880 3.580 4.220 5.280 ;
        RECT  2.490 3.360 2.830 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.740 1.180 3.050 1.410 ;
        RECT  0.740 1.180 1.080 1.520 ;
        RECT  2.060 1.180 3.050 1.520 ;
        RECT  2.820 2.015 3.350 2.355 ;
        RECT  2.820 1.180 3.050 3.130 ;
        RECT  1.330 2.900 3.050 3.130 ;
        RECT  1.330 2.900 1.670 3.960 ;
        RECT  0.740 1.180 2.90 1.410 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.823  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 1.230 2.565 2.980 ;
        RECT  2.000 2.690 2.400 3.240 ;
        RECT  2.070 1.230 2.565 1.570 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.805 2.205 1.310 2.630 ;
        RECT  0.995 1.870 1.310 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.105 0.575 2.460 ;
        RECT  0.125 1.640 0.505 2.460 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 0.710 ;
        RECT  1.300 -0.400 1.640 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.630 3.265 2.970 5.280 ;
        RECT  1.330 3.320 1.670 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.740 1.205 1.770 1.545 ;
        RECT  1.540 2.015 2.100 2.355 ;
        RECT  1.540 1.205 1.770 3.090 ;
        RECT  0.180 2.860 1.770 3.090 ;
        RECT  0.180 2.860 0.520 3.960 ;
    END
END OR2X2

MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.770  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.860 2.405 3.390 ;
        RECT  2.175 1.115 2.405 3.390 ;
        RECT  2.000 1.115 2.405 1.455 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.905 1.600 1.290 2.230 ;
        RECT  0.755 1.600 1.290 2.020 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.195 0.605 2.695 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  1.095 -0.400 1.435 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  1.370 3.610 1.710 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.025 1.750 1.365 ;
        RECT  1.520 2.015 1.945 2.355 ;
        RECT  1.520 1.025 1.750 3.325 ;
        RECT  0.180 3.095 1.750 3.325 ;
        RECT  0.180 3.095 0.520 3.520 ;
    END
END OR2X1

MACRO OR2X0
    CLASS CORE ;
    FOREIGN OR2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.558  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.860 2.405 3.390 ;
        RECT  2.175 0.630 2.405 3.390 ;
        RECT  2.000 0.630 2.405 0.970 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.195 0.605 2.690 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.905 1.600 1.290 2.230 ;
        RECT  0.755 1.600 1.290 2.020 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  1.200 3.690 1.540 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.665 1.025 1.750 1.365 ;
        RECT  1.520 2.015 1.945 2.355 ;
        RECT  1.520 1.025 1.750 3.325 ;
        RECT  0.370 3.095 1.750 3.325 ;
        RECT  0.370 3.095 0.710 4.030 ;
    END
END OR2X0

MACRO ON33X4
    CLASS CORE ;
    FOREIGN ON33X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.100 4.285 2.710 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.655 3.240 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.050 3.045 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 2.110 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 0.780 8.065 3.960 ;
        RECT  6.390 2.050 8.065 2.280 ;
        RECT  6.230 2.640 6.620 3.750 ;
        RECT  6.390 1.110 6.620 3.750 ;
        RECT  6.230 1.110 6.620 1.450 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.950 -0.400 7.290 1.700 ;
        RECT  5.680 -0.400 6.020 0.710 ;
        RECT  1.540 -0.400 1.880 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.950 2.640 7.290 5.280 ;
        RECT  5.670 4.160 6.010 5.280 ;
        RECT  4.210 3.930 4.550 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.920 1.700 ;
        RECT  2.900 0.790 4.735 1.130 ;
        RECT  4.505 0.790 4.735 1.960 ;
        RECT  4.515 1.930 4.990 2.270 ;
        RECT  4.515 1.770 4.745 3.190 ;
        RECT  3.885 2.960 4.745 3.190 ;
        RECT  3.885 2.960 4.115 3.700 ;
        RECT  2.335 3.470 4.115 3.700 ;
        RECT  2.335 2.860 2.675 4.140 ;
        RECT  4.965 1.360 5.450 1.700 ;
        RECT  5.220 1.945 6.160 2.285 ;
        RECT  5.220 1.360 5.450 3.585 ;
        RECT  4.910 3.355 5.250 4.180 ;
        RECT  0.860 1.360 2.40 1.700 ;
    END
END ON33X4

MACRO ON33X2
    CLASS CORE ;
    FOREIGN ON33X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.090 3.470 3.430 3.880 ;
        RECT  2.645 3.470 3.430 3.850 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.910 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 3.470 4.580 3.880 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 5.180 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.155 3.460 5.740 3.890 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.120 6.355 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.640 1.135 3.560 ;
        RECT  0.740 1.250 1.080 1.590 ;
        RECT  0.740 1.250 0.970 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.430 6.750 5.280 ;
        RECT  2.570 4.080 2.910 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  2.770 -0.400 4.230 0.950 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.960 1.250 2.400 1.590 ;
        RECT  1.200 2.070 2.190 2.410 ;
        RECT  1.960 1.250 2.190 3.560 ;
        RECT  1.960 2.640 2.400 3.560 ;
        RECT  4.590 0.630 4.930 1.700 ;
        RECT  3.330 1.360 6.190 1.700 ;
        RECT  5.290 0.630 6.815 0.950 ;
        RECT  2.420 2.070 2.870 2.410 ;
        RECT  2.630 2.070 2.870 3.200 ;
        RECT  6.585 0.630 6.815 3.200 ;
        RECT  2.630 2.860 6.815 3.200 ;
        RECT  3.330 1.360 5.60 1.700 ;
        RECT  2.630 2.860 5.50 3.200 ;
    END
END ON33X2

MACRO ON33X1
    CLASS CORE ;
    FOREIGN ON33X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.040 3.655 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.035 4.305 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.911  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 2.860 4.915 3.240 ;
        RECT  4.535 0.790 4.915 3.240 ;
        RECT  4.300 0.790 4.915 1.700 ;
        RECT  2.900 0.790 4.915 1.130 ;
        RECT  2.335 2.860 2.675 4.140 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.285 2.860 1.765 3.240 ;
        RECT  1.285 2.120 1.625 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.935 2.060 2.395 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.060 3.045 2.630 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.540 -0.400 1.880 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.355 3.515 4.695 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.920 1.700 ;
        RECT  0.860 1.360 2.30 1.700 ;
    END
END ON33X1

MACRO ON33X0
    CLASS CORE ;
    FOREIGN ON33X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.855 1.155 3.240 ;
        RECT  0.835 2.240 1.155 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.255 1.925 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.860 2.630 3.260 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.620 2.155 3.185 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.135 2.860 3.675 3.260 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.840 3.510 4.235 3.850 ;
        RECT  3.905 0.630 4.235 3.850 ;
        RECT  2.520 0.630 4.235 0.950 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.505 3.010 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.505 4.080 3.845 5.280 ;
        RECT  0.220 3.545 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.120 -0.400 1.460 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.820 0.630 2.160 1.590 ;
        RECT  0.445 1.220 2.160 1.590 ;
        RECT  0.445 1.250 3.460 1.590 ;
        RECT  0.445 1.250 2.40 1.590 ;
    END
END ON33X0

MACRO ON333X1
    CLASS CORE ;
    FOREIGN ON333X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.070 5.565 2.680 ;
        END
    END H
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.744  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 3.470 6.805 3.755 ;
        RECT  6.540 1.360 6.805 3.755 ;
        RECT  6.280 2.860 6.805 3.755 ;
        RECT  4.995 1.360 6.805 1.700 ;
        RECT  2.335 2.860 2.675 4.140 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 4.935 3.240 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.115 4.305 2.695 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.655 3.240 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.060 3.045 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.920 2.110 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.120 6.310 2.630 ;
        END
    END J
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.330 3.985 4.670 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  1.540 -0.400 1.880 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.920 1.700 ;
        RECT  2.900 0.790 6.070 1.130 ;
        RECT  0.860 1.360 2.60 1.700 ;
        RECT  2.900 0.790 5.50 1.130 ;
    END
END ON333X1

MACRO ON333X0
    CLASS CORE ;
    FOREIGN ON333X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.555 1.850 1.975 2.190 ;
        RECT  1.385 3.460 1.785 3.850 ;
        RECT  1.555 1.850 1.785 3.850 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.860 2.775 3.260 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.930 1.970 3.310 2.310 ;
        RECT  2.645 2.250 3.160 2.630 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.930 2.250 1.270 2.780 ;
        RECT  0.755 2.250 1.270 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.270 2.860 3.885 3.265 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.640 2.460 ;
        RECT  3.905 2.120 4.285 2.630 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.282  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.155 3.555 6.185 3.895 ;
        RECT  5.955 0.710 6.185 3.895 ;
        RECT  5.795 3.470 6.185 3.895 ;
        RECT  4.550 0.710 6.185 1.030 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.530 2.855 5.115 3.270 ;
        END
    END H
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.440 2.250 5.725 2.890 ;
        RECT  5.165 2.250 5.725 2.630 ;
        END
    END J
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.685 0.525 3.280 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.250 -0.400 1.590 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  3.820 4.125 4.160 5.280 ;
        RECT  0.535 3.570 0.875 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.650 1.170 2.290 1.410 ;
        RECT  1.950 0.710 2.290 1.410 ;
        RECT  0.650 1.170 0.990 1.510 ;
        RECT  1.995 1.330 3.590 1.615 ;
        RECT  3.250 1.330 3.590 1.670 ;
        RECT  2.650 0.710 4.195 1.030 ;
        RECT  3.965 0.710 4.195 1.600 ;
        RECT  3.965 1.260 5.590 1.600 ;
    END
END ON333X0

MACRO ON332X1
    CLASS CORE ;
    FOREIGN ON332X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.935 2.100 2.395 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.060 3.045 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.655 3.240 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.115 4.305 2.695 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 4.935 3.240 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 3.470 6.175 3.755 ;
        RECT  5.910 1.360 6.175 3.755 ;
        RECT  5.650 2.860 6.175 3.755 ;
        RECT  5.020 1.360 6.175 1.700 ;
        RECT  2.335 2.860 2.675 4.140 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.120 5.680 2.630 ;
        END
    END H
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.540 -0.400 1.880 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.355 3.985 4.695 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.920 1.700 ;
        RECT  2.900 0.790 6.120 1.130 ;
        RECT  0.860 1.360 2.20 1.700 ;
        RECT  2.900 0.790 5.60 1.130 ;
    END
END ON332X1

MACRO ON332X0
    CLASS CORE ;
    FOREIGN ON332X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.835 2.230 1.230 2.780 ;
        RECT  0.755 2.230 1.230 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.485 1.770 1.905 2.110 ;
        RECT  1.385 3.460 1.715 3.850 ;
        RECT  1.485 1.770 1.715 3.850 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.855 2.595 3.275 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.970 3.190 2.315 ;
        RECT  2.645 1.970 3.025 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.230 2.850 3.760 3.275 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.200 4.485 2.630 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.959  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 3.550 5.545 3.890 ;
        RECT  5.315 1.130 5.545 3.890 ;
        RECT  5.165 3.470 5.545 3.890 ;
        RECT  4.525 1.130 5.545 1.470 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.855 5.060 3.265 ;
        END
    END H
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.770 0.570 3.290 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  1.125 -0.400 1.465 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.625 4.170 3.965 5.280 ;
        RECT  0.220 3.570 0.560 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.170 2.165 1.410 ;
        RECT  1.825 0.630 2.165 1.410 ;
        RECT  0.445 1.170 0.785 1.510 ;
        RECT  1.975 1.250 3.465 1.535 ;
        RECT  3.125 1.250 3.465 1.590 ;
        RECT  2.525 0.630 4.065 0.950 ;
    END
END ON332X0

MACRO ON331X1
    CLASS CORE ;
    FOREIGN ON331X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 3.470 5.545 3.755 ;
        RECT  5.150 0.885 5.545 3.755 ;
        RECT  4.980 0.885 5.545 1.700 ;
        RECT  2.335 2.860 2.675 4.140 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 4.920 3.240 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.115 4.305 2.695 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.655 3.240 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.060 3.045 2.630 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.935 2.100 2.395 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.355 3.985 4.695 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  1.540 -0.400 1.880 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.920 1.700 ;
        RECT  0.860 1.360 2.40 1.700 ;
        RECT  2.900 0.790 4.600 1.130 ;
    END
END ON331X1

MACRO ON331X0
    CLASS CORE ;
    FOREIGN ON331X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.135 3.850 ;
        RECT  0.795 2.300 1.135 3.850 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.195 1.935 2.635 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.855 2.595 3.270 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.970 3.160 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.160 2.860 3.680 3.265 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.165 4.355 2.640 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.840 3.520 4.915 3.860 ;
        RECT  4.585 1.170 4.915 3.860 ;
        RECT  4.535 3.470 4.915 3.860 ;
        RECT  4.520 1.170 4.915 1.510 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.715 0.505 3.250 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.120 -0.400 1.460 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.505 4.120 3.845 5.280 ;
        RECT  0.220 3.570 0.525 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.820 0.630 2.160 1.590 ;
        RECT  0.445 1.170 2.160 1.590 ;
        RECT  0.445 1.250 3.460 1.590 ;
        RECT  2.520 0.630 4.075 0.950 ;
        RECT  0.445 1.250 2.80 1.590 ;
    END
END ON331X0

MACRO ON32X4
    CLASS CORE ;
    FOREIGN ON32X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.030 3.655 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.455  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.050 3.045 2.630 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 2.110 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 0.780 7.435 3.960 ;
        RECT  5.760 2.050 7.435 2.280 ;
        RECT  5.600 2.640 5.990 3.750 ;
        RECT  5.760 1.110 5.990 3.750 ;
        RECT  5.600 1.110 5.990 1.450 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.700 ;
        RECT  5.050 -0.400 5.390 0.710 ;
        RECT  1.540 -0.400 1.880 1.160 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 2.640 6.660 5.280 ;
        RECT  5.040 4.160 5.380 5.280 ;
        RECT  3.540 3.320 3.880 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.620 0.740 3.960 1.080 ;
        RECT  2.220 0.850 3.960 1.080 ;
        RECT  0.860 1.360 1.200 1.700 ;
        RECT  2.220 0.850 2.560 1.700 ;
        RECT  0.860 1.470 2.560 1.700 ;
        RECT  2.940 1.360 3.280 1.700 ;
        RECT  2.940 1.470 4.105 1.700 ;
        RECT  3.875 1.470 4.105 1.960 ;
        RECT  3.885 1.930 4.360 2.270 ;
        RECT  3.885 1.770 4.115 3.090 ;
        RECT  2.335 2.860 4.115 3.090 ;
        RECT  2.335 2.860 2.675 4.020 ;
        RECT  4.335 1.360 4.820 1.700 ;
        RECT  4.590 1.945 5.530 2.285 ;
        RECT  4.590 1.360 4.820 3.585 ;
        RECT  4.280 3.355 4.620 4.180 ;
    END
END ON32X4

MACRO ON32X2
    CLASS CORE ;
    FOREIGN ON32X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.090 3.470 3.430 3.880 ;
        RECT  2.645 3.470 3.430 3.850 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.845 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 3.470 4.530 3.880 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.160 3.415 5.680 3.885 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.640 1.135 3.560 ;
        RECT  0.740 1.250 1.080 1.590 ;
        RECT  0.740 1.250 0.970 3.560 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 5.080 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.910 2.790 6.140 5.280 ;
        RECT  5.650 2.790 6.140 3.130 ;
        RECT  2.570 4.080 2.910 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  3.890 -0.400 4.230 0.950 ;
        RECT  2.610 1.350 2.950 1.690 ;
        RECT  2.670 -0.400 2.950 1.690 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.960 0.640 2.440 0.980 ;
        RECT  1.200 2.070 2.190 2.410 ;
        RECT  1.960 0.640 2.190 3.560 ;
        RECT  1.960 2.640 2.400 3.560 ;
        RECT  5.150 1.350 5.490 1.870 ;
        RECT  4.075 1.640 5.490 1.870 ;
        RECT  2.420 2.070 2.870 2.410 ;
        RECT  2.630 2.070 2.870 3.200 ;
        RECT  4.075 1.640 4.305 3.200 ;
        RECT  2.630 2.860 4.770 3.200 ;
        RECT  4.590 0.630 6.050 0.950 ;
        RECT  3.190 0.630 3.530 1.410 ;
        RECT  4.590 0.630 4.870 1.410 ;
        RECT  3.190 1.180 4.870 1.410 ;
        RECT  2.630 2.860 3.80 3.200 ;
    END
END ON32X2

MACRO ON32X1
    CLASS CORE ;
    FOREIGN ON32X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.860 1.480 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 2.860 2.395 3.240 ;
        RECT  1.860 2.120 2.200 3.240 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.570 2.110 3.035 2.640 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.655 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.340  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.250 4.285 2.630 ;
        RECT  2.120 3.475 4.125 3.760 ;
        RECT  3.895 1.480 4.125 3.760 ;
        RECT  3.060 1.480 4.125 1.710 ;
        RECT  3.060 1.360 3.400 1.710 ;
        RECT  2.120 3.475 2.460 3.815 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.765 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.530 3.990 3.870 5.280 ;
        RECT  0.180 3.100 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.620 -0.400 1.960 1.250 ;
        RECT  0.180 -0.400 0.520 1.250 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.340 0.900 4.120 1.130 ;
        RECT  3.780 0.900 4.120 1.250 ;
        RECT  0.900 1.360 1.240 1.710 ;
        RECT  2.340 0.900 2.680 1.710 ;
        RECT  0.900 1.480 2.680 1.710 ;
    END
END ON32X1

MACRO ON32X0
    CLASS CORE ;
    FOREIGN ON32X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.155 3.850 ;
        RECT  0.835 2.580 1.155 3.850 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.195 1.935 2.635 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.181  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.860 2.605 3.270 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.181  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.170 3.170 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.742  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.840 3.595 3.655 3.935 ;
        RECT  3.400 1.210 3.655 3.935 ;
        RECT  3.265 3.470 3.655 3.935 ;
        RECT  2.520 1.210 3.655 1.550 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.860 0.505 3.410 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.070 4.170 3.410 5.280 ;
        RECT  0.185 3.670 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  1.120 -0.400 1.460 0.790 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.820 0.710 2.160 1.590 ;
        RECT  0.445 1.250 2.160 1.590 ;
    END
END ON32X0

MACRO ON322X1
    CLASS CORE ;
    FOREIGN ON322X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 2.105 2.410 2.645 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.205 2.115 3.675 2.635 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.285 3.240 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.115 4.935 2.695 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.120 5.610 2.460 ;
        RECT  5.165 2.120 5.555 3.240 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.632  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.200 3.475 6.175 3.760 ;
        RECT  5.785 2.860 6.175 3.760 ;
        RECT  5.840 1.390 6.070 3.760 ;
        RECT  4.890 1.390 6.070 1.620 ;
        RECT  5.780 3.335 6.175 3.760 ;
        RECT  4.890 1.280 5.230 1.620 ;
        RECT  2.970 2.895 3.310 3.760 ;
        RECT  2.200 2.895 2.540 3.760 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.540 -0.400 1.880 1.160 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.320 3.990 4.660 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 1.200 1.700 ;
        RECT  2.220 1.360 2.560 1.700 ;
        RECT  3.530 1.360 3.880 1.700 ;
        RECT  0.860 1.470 3.880 1.700 ;
        RECT  2.845 0.740 5.910 0.970 ;
        RECT  2.845 0.740 3.185 1.080 ;
        RECT  4.205 0.740 4.550 1.080 ;
        RECT  5.570 0.740 5.910 1.080 ;
        RECT  0.860 1.470 2.70 1.700 ;
        RECT  2.845 0.740 4.00 0.970 ;
    END
END ON322X1

MACRO ON322X0
    CLASS CORE ;
    FOREIGN ON322X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.220 1.345 2.640 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.920 1.905 3.260 ;
        RECT  1.385 2.920 1.775 3.850 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.585 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.860 3.260 3.280 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 2.190 3.825 2.630 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.955  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 3.550 4.915 3.890 ;
        RECT  4.685 1.130 4.915 3.890 ;
        RECT  4.535 3.470 4.915 3.890 ;
        RECT  4.025 1.130 4.915 1.470 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.850 4.430 3.260 ;
        END
    END G
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.770 0.565 3.290 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.125 -0.400 1.465 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.195 4.125 3.535 5.280 ;
        RECT  0.220 3.570 0.560 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.825 0.630 2.165 1.510 ;
        RECT  0.445 1.170 2.165 1.510 ;
        RECT  2.525 0.630 3.680 0.950 ;
        RECT  2.525 0.630 2.865 1.740 ;
    END
END ON322X0

MACRO ON321X4
    CLASS CORE ;
    FOREIGN ON321X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.900 2.105 2.410 2.645 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.080 3.385 2.635 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.435  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.770 2.120 4.285 3.240 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.020 4.905 2.630 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.100 2.860 1.765 3.240 ;
        RECT  1.100 2.120 1.440 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 0.780 8.695 3.960 ;
        RECT  7.020 2.050 8.695 2.280 ;
        RECT  6.860 2.640 7.250 3.750 ;
        RECT  7.020 1.110 7.250 3.750 ;
        RECT  6.860 1.110 7.250 1.450 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 2.640 7.920 5.280 ;
        RECT  6.300 4.160 6.640 5.280 ;
        RECT  4.045 3.990 4.385 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.700 ;
        RECT  6.310 -0.400 6.650 0.710 ;
        RECT  1.540 -0.400 1.880 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.880 1.700 ;
        RECT  2.845 0.740 4.550 1.080 ;
        RECT  4.930 0.740 5.365 1.080 ;
        RECT  5.135 1.930 5.620 2.270 ;
        RECT  5.135 0.740 5.365 3.090 ;
        RECT  2.345 2.895 2.685 3.760 ;
        RECT  4.840 2.860 5.180 3.760 ;
        RECT  2.345 3.475 5.180 3.760 ;
        RECT  5.595 1.360 6.080 1.700 ;
        RECT  5.850 1.945 6.790 2.285 ;
        RECT  5.850 1.360 6.080 3.520 ;
        RECT  5.540 3.290 5.880 4.180 ;
        RECT  0.860 1.360 2.60 1.700 ;
        RECT  2.345 3.475 4.50 3.760 ;
    END
END ON321X4

MACRO ON321X2
    CLASS CORE ;
    FOREIGN ON321X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.785 2.120 4.285 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.390 3.430 4.925 3.890 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.920 2.080 5.545 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.050 6.195 2.630 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.450 3.655 4.090 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.750 1.135 3.560 ;
        RECT  0.740 1.250 1.080 1.590 ;
        RECT  0.740 1.250 0.970 3.560 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.080 6.920 2.630 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.870 3.320 6.680 5.280 ;
        RECT  2.760 2.860 3.095 3.200 ;
        RECT  2.760 2.860 3.045 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  2.760 -0.400 4.220 0.950 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.940 1.250 2.400 1.590 ;
        RECT  1.200 1.945 2.170 2.285 ;
        RECT  1.940 1.250 2.170 3.560 ;
        RECT  1.940 2.750 2.400 3.560 ;
        RECT  3.320 1.360 6.300 1.700 ;
        RECT  5.400 0.630 7.110 0.950 ;
        RECT  6.770 1.330 7.380 1.670 ;
        RECT  2.410 1.945 3.555 2.285 ;
        RECT  3.325 1.945 3.555 3.090 ;
        RECT  3.325 2.860 7.380 3.090 ;
        RECT  4.650 2.860 4.990 3.200 ;
        RECT  7.150 1.330 7.380 3.780 ;
        RECT  7.040 2.860 7.380 3.780 ;
        RECT  3.320 1.360 5.60 1.700 ;
        RECT  3.325 2.860 6.60 3.090 ;
    END
END ON321X2

MACRO ON321X1
    CLASS CORE ;
    FOREIGN ON321X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.760 2.120 2.395 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.810 3.045 3.240 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.080 3.675 2.690 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.369  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.455 2.460 ;
        RECT  3.905 1.640 4.285 2.460 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.976  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 2.690 4.925 3.875 ;
        RECT  4.685 1.290 4.925 3.875 ;
        RECT  4.520 1.290 4.925 1.630 ;
        RECT  2.055 3.515 4.925 3.795 ;
        RECT  4.515 2.690 4.925 3.795 ;
        RECT  2.055 2.860 2.395 3.910 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.090 2.860 1.765 3.240 ;
        RECT  1.090 2.120 1.430 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.575 4.025 3.915 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.415 -0.400 1.755 1.040 ;
        RECT  0.180 -0.400 0.520 1.040 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.800 1.290 3.640 1.580 ;
        RECT  0.800 1.290 2.370 1.630 ;
        RECT  3.290 1.290 3.640 1.630 ;
        RECT  2.675 0.700 4.245 1.040 ;
        RECT  0.800 1.290 2.30 1.580 ;
    END
END ON321X1

MACRO ON321X0
    CLASS CORE ;
    FOREIGN ON321X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.680 1.640 1.135 2.160 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.075 1.840 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.860 2.605 3.240 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.170 3.170 2.630 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.155  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.860 3.750 3.240 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.857  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.800 3.490 4.285 3.830 ;
        RECT  3.980 0.630 4.285 3.830 ;
        RECT  3.615 0.630 4.285 0.950 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.795 0.600 3.300 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  2.990 4.070 3.330 5.280 ;
        RECT  0.220 3.570 0.560 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.185 -0.400 1.525 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.885 0.630 2.225 1.410 ;
        RECT  0.490 1.070 2.225 1.410 ;
        RECT  0.490 1.180 3.485 1.410 ;
        RECT  3.145 1.180 3.485 1.810 ;
        RECT  0.490 1.180 2.20 1.410 ;
    END
END ON321X0

MACRO ON31X4
    CLASS CORE ;
    FOREIGN ON31X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.070 3.025 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 2.110 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 0.780 6.805 3.960 ;
        RECT  5.130 2.050 6.805 2.280 ;
        RECT  4.970 2.640 5.360 3.750 ;
        RECT  5.130 1.110 5.360 3.750 ;
        RECT  4.970 1.110 5.360 1.450 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.700 ;
        RECT  4.420 -0.400 4.760 0.710 ;
        RECT  1.540 -0.400 1.880 1.160 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 2.640 6.030 5.280 ;
        RECT  4.410 4.160 4.750 5.280 ;
        RECT  2.950 3.320 3.290 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 1.200 1.700 ;
        RECT  2.220 1.360 2.560 1.700 ;
        RECT  0.860 1.470 2.560 1.700 ;
        RECT  2.940 0.740 3.280 1.700 ;
        RECT  3.245 1.470 3.475 2.000 ;
        RECT  3.255 1.930 3.730 2.270 ;
        RECT  3.255 1.930 3.485 3.090 ;
        RECT  2.150 2.860 3.485 3.090 ;
        RECT  2.150 2.860 2.490 4.180 ;
        RECT  3.650 0.780 4.190 1.120 ;
        RECT  3.705 0.780 4.190 1.700 ;
        RECT  3.960 1.945 4.900 2.285 ;
        RECT  3.960 0.780 4.190 3.485 ;
        RECT  3.650 3.255 3.990 4.180 ;
    END
END ON31X4

MACRO ON31X2
    CLASS CORE ;
    FOREIGN ON31X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.090 3.470 3.430 3.880 ;
        RECT  2.645 3.470 3.430 3.850 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.845 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 3.470 4.530 3.880 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 5.180 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.640 1.135 3.560 ;
        RECT  0.740 1.250 1.080 1.590 ;
        RECT  0.740 1.250 0.970 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 2.860 5.490 5.280 ;
        RECT  2.570 4.080 2.910 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.890 -0.400 4.230 0.950 ;
        RECT  2.610 1.350 2.950 1.690 ;
        RECT  2.670 -0.400 2.950 1.690 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.960 0.640 2.440 0.980 ;
        RECT  1.200 2.070 2.190 2.410 ;
        RECT  1.960 0.640 2.190 3.560 ;
        RECT  1.960 2.640 2.400 3.560 ;
        RECT  4.590 0.630 4.930 0.950 ;
        RECT  3.190 0.630 3.530 1.410 ;
        RECT  4.590 0.630 4.920 1.410 ;
        RECT  3.190 1.180 4.920 1.410 ;
        RECT  5.150 1.350 5.490 1.870 ;
        RECT  4.075 1.640 5.490 1.870 ;
        RECT  2.420 2.070 2.870 2.410 ;
        RECT  2.630 2.070 2.870 3.200 ;
        RECT  4.075 1.640 4.305 3.200 ;
        RECT  2.630 2.860 4.770 3.200 ;
        RECT  2.630 2.860 3.40 3.200 ;
    END
END ON31X2

MACRO ON31X1
    CLASS CORE ;
    FOREIGN ON31X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.860 1.480 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 2.120 2.395 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.120 3.025 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.338  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.655 2.630 ;
        RECT  2.120 3.475 3.605 3.705 ;
        RECT  3.275 1.360 3.605 3.705 ;
        RECT  3.060 1.360 3.605 1.710 ;
        RECT  2.120 3.475 2.460 4.180 ;
        RECT  2.120 3.370 2.455 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.765 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.920 3.990 3.260 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  1.620 -0.400 1.960 1.250 ;
        RECT  0.180 -0.400 0.520 1.475 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.360 1.240 1.710 ;
        RECT  2.340 0.900 2.680 1.710 ;
        RECT  0.900 1.480 2.680 1.710 ;
    END
END ON31X1

MACRO ON31X0
    CLASS CORE ;
    FOREIGN ON31X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.135 2.185 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.805 1.835 2.145 ;
        RECT  1.385 1.805 1.780 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.142  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.440 2.500 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.622  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.640 3.470 3.025 3.860 ;
        RECT  2.730 1.285 3.025 3.860 ;
        RECT  2.630 1.285 3.025 1.625 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.194  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.370 0.505 3.290 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.440 4.170 2.780 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.155 -0.400 1.495 0.745 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.855 0.670 2.195 1.355 ;
        RECT  0.525 1.015 2.195 1.355 ;
    END
END ON31X0

MACRO ON311X4
    CLASS CORE ;
    FOREIGN ON311X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 2.120 2.395 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.270 1.980 3.645 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.000 3.040 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.860 1.765 3.240 ;
        RECT  1.140 2.120 1.480 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 0.780 7.435 3.960 ;
        RECT  5.760 2.050 7.435 2.280 ;
        RECT  5.600 2.640 5.990 3.750 ;
        RECT  5.760 1.110 5.990 3.750 ;
        RECT  5.600 1.110 5.990 1.450 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 2.640 6.660 5.280 ;
        RECT  5.040 4.160 5.380 5.280 ;
        RECT  2.905 3.320 3.245 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.700 ;
        RECT  5.050 -0.400 5.390 0.710 ;
        RECT  1.620 -0.400 1.960 1.240 ;
        RECT  0.180 -0.400 0.520 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 0.820 1.240 1.700 ;
        RECT  2.340 0.820 2.680 1.700 ;
        RECT  0.900 1.470 2.680 1.700 ;
        RECT  3.535 0.820 4.105 1.700 ;
        RECT  3.875 1.930 4.360 2.270 ;
        RECT  2.105 2.860 4.105 3.090 ;
        RECT  3.875 0.820 4.105 3.195 ;
        RECT  3.665 2.860 4.105 3.195 ;
        RECT  2.105 2.860 2.445 4.180 ;
        RECT  4.335 0.780 4.820 1.700 ;
        RECT  4.590 1.945 5.530 2.285 ;
        RECT  4.590 0.780 4.820 3.600 ;
        RECT  4.280 3.370 4.620 4.180 ;
        RECT  2.105 2.860 3.80 3.090 ;
    END
END ON311X4

MACRO ON311X2
    CLASS CORE ;
    FOREIGN ON311X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.605 2.120 4.285 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.280 3.430 4.905 3.880 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.120 6.185 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.120 5.545 2.630 ;
        RECT  4.975 2.120 5.545 2.460 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.205 3.450 3.655 4.090 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.640 1.135 3.560 ;
        RECT  0.740 1.250 1.080 1.590 ;
        RECT  0.740 1.250 0.970 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.135 3.440 5.420 5.280 ;
        RECT  2.635 3.300 2.975 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  2.760 -0.400 4.220 0.950 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.940 1.250 2.400 1.590 ;
        RECT  1.200 2.070 2.170 2.410 ;
        RECT  1.940 1.250 2.170 2.980 ;
        RECT  1.940 2.640 2.400 2.980 ;
        RECT  4.615 0.630 4.955 1.410 ;
        RECT  3.320 1.180 4.955 1.410 ;
        RECT  3.320 1.180 3.660 1.700 ;
        RECT  5.780 1.360 6.120 1.890 ;
        RECT  4.515 1.660 6.120 1.890 ;
        RECT  2.410 2.070 3.375 2.410 ;
        RECT  4.515 1.660 4.745 3.090 ;
        RECT  3.145 2.070 3.375 3.090 ;
        RECT  4.515 2.700 4.860 3.090 ;
        RECT  3.145 2.860 6.120 3.090 ;
        RECT  5.780 2.860 6.120 3.780 ;
        RECT  3.145 2.860 5.40 3.090 ;
    END
END ON311X2

MACRO ON311X1
    CLASS CORE ;
    FOREIGN ON311X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.380 2.630 ;
        RECT  1.040 1.845 1.380 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.610 2.010 2.055 2.350 ;
        RECT  1.385 2.860 1.875 3.240 ;
        RECT  1.610 2.010 1.875 3.240 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.374  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.385 2.100 3.025 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.374  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.470 3.655 4.250 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.648  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.115 2.970 3.645 3.220 ;
        RECT  3.255 1.320 3.645 3.220 ;
        RECT  3.250 2.880 3.645 3.220 ;
        RECT  3.250 1.320 3.645 1.660 ;
        RECT  1.895 3.470 2.395 3.850 ;
        RECT  2.115 2.970 2.395 3.850 ;
        RECT  1.925 3.465 2.395 3.850 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.505 2.460 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.480 4.170 2.835 5.280 ;
        RECT  0.180 2.900 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  1.420 -0.400 1.760 1.040 ;
        RECT  0.180 -0.400 0.520 1.040 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.800 1.320 2.440 1.610 ;
        RECT  0.800 1.320 1.140 1.615 ;
        RECT  2.100 1.320 2.440 1.660 ;
    END
END ON311X1

MACRO ON311X0
    CLASS CORE ;
    FOREIGN ON311X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.975 1.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.580 1.765 3.240 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.155  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.095 2.510 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.155  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.215 3.650 2.810 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.836  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.740 3.420 3.580 3.750 ;
        RECT  2.740 1.170 3.500 1.510 ;
        RECT  1.640 3.470 3.025 3.850 ;
        RECT  2.740 1.170 2.990 3.850 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.207  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.610 0.505 3.240 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.440 4.090 2.780 5.280 ;
        RECT  0.180 4.105 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  1.185 -0.400 1.525 0.835 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.170 2.260 1.510 ;
    END
END ON311X0

MACRO ON22X4
    CLASS CORE ;
    FOREIGN ON22X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.100 0.670 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.100 3.160 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.050 2.415 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.360 2.040 1.765 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 0.780 6.805 3.960 ;
        RECT  5.130 2.050 6.805 2.280 ;
        RECT  4.970 2.640 5.360 3.750 ;
        RECT  5.130 1.110 5.360 3.750 ;
        RECT  4.970 1.110 5.360 1.450 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 2.640 6.030 5.280 ;
        RECT  4.410 4.160 4.750 5.280 ;
        RECT  2.950 3.350 3.290 5.280 ;
        RECT  0.420 3.320 0.760 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.700 ;
        RECT  4.420 -0.400 4.760 0.710 ;
        RECT  2.340 -0.400 2.680 1.200 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.820 1.960 1.050 ;
        RECT  1.620 0.820 1.960 1.660 ;
        RECT  0.180 0.820 0.520 1.660 ;
        RECT  3.060 0.820 3.400 1.660 ;
        RECT  1.620 1.430 3.400 1.660 ;
        RECT  0.900 1.280 1.240 1.620 ;
        RECT  3.730 2.120 4.070 2.460 ;
        RECT  0.900 1.280 1.130 3.090 ;
        RECT  3.730 2.120 3.960 3.090 ;
        RECT  0.900 2.860 3.960 3.090 ;
        RECT  1.720 2.860 2.060 4.140 ;
        RECT  3.650 1.360 4.530 1.700 ;
        RECT  4.300 1.945 4.900 2.285 ;
        RECT  4.300 1.360 4.530 3.585 ;
        RECT  3.650 3.355 4.530 3.585 ;
        RECT  3.650 3.355 3.990 4.180 ;
        RECT  0.900 2.860 2.90 3.090 ;
    END
END ON22X4

MACRO ON22X2
    CLASS CORE ;
    FOREIGN ON22X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 2.250 3.705 2.760 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.640 1.240 3.560 ;
        RECT  0.755 1.250 1.240 1.590 ;
        RECT  0.755 1.250 0.985 3.560 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.460 2.120 6.175 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 5.075 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.875 3.460 4.350 3.980 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.215 -0.400 5.555 1.530 ;
        RECT  1.620 -0.400 1.960 1.560 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.645 2.995 5.985 5.280 ;
        RECT  3.070 2.990 3.415 5.280 ;
        RECT  1.620 2.640 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.190 1.255 2.680 1.595 ;
        RECT  1.380 1.945 2.420 2.285 ;
        RECT  2.190 1.255 2.420 3.560 ;
        RECT  2.190 2.640 2.680 3.560 ;
        RECT  2.805 1.790 4.235 2.020 ;
        RECT  3.895 1.190 4.235 2.020 ;
        RECT  2.650 1.945 3.035 2.285 ;
        RECT  3.935 1.190 4.235 3.200 ;
        RECT  3.935 2.860 4.565 3.200 ;
    END
END ON22X2

MACRO ON22X1
    CLASS CORE ;
    FOREIGN ON22X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 2.065 1.780 2.675 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.405 3.240 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.080 3.080 2.660 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.920 3.475 1.960 3.815 ;
        RECT  0.900 1.360 1.240 1.700 ;
        RECT  0.920 1.360 1.150 3.815 ;
        RECT  0.755 2.860 1.150 3.240 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.690 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.015 3.010 3.355 5.280 ;
        RECT  0.180 3.100 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.340 -0.400 2.680 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.900 1.970 1.130 ;
        RECT  0.180 0.900 0.520 1.520 ;
        RECT  1.620 0.900 1.970 1.800 ;
        RECT  3.060 1.180 3.400 1.800 ;
        RECT  1.620 1.570 3.400 1.800 ;
    END
END ON22X1

MACRO ON22X0
    CLASS CORE ;
    FOREIGN ON22X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.490 0.505 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 2.195 1.305 2.635 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.855 1.935 3.260 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.030 3.025 2.645 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.649  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 3.620 2.395 3.960 ;
        RECT  2.165 1.780 2.395 3.960 ;
        RECT  2.015 3.520 2.395 3.960 ;
        RECT  2.020 3.475 2.395 3.960 ;
        RECT  1.525 1.780 2.395 2.010 ;
        RECT  1.525 1.210 1.755 2.010 ;
        RECT  0.625 1.210 1.755 1.550 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.625 3.620 2.910 5.280 ;
        RECT  0.220 3.620 0.560 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.030 -0.400 2.370 1.550 ;
        END
    END gnd!
END ON22X0

MACRO ON222X4
    CLASS CORE ;
    FOREIGN ON222X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.340 2.120 1.765 3.240 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.780 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.160 2.120 3.675 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.285 3.240 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.060 4.905 2.680 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.960 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 0.780 8.695 3.960 ;
        RECT  7.020 2.050 8.695 2.280 ;
        RECT  6.860 2.640 7.250 3.750 ;
        RECT  7.020 1.110 7.250 3.750 ;
        RECT  6.860 1.110 7.250 1.450 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 2.640 7.920 5.280 ;
        RECT  6.300 4.160 6.640 5.280 ;
        RECT  3.535 3.930 3.875 5.280 ;
        RECT  0.375 2.860 0.715 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.700 ;
        RECT  6.310 -0.400 6.650 0.710 ;
        RECT  1.540 -0.400 1.880 1.125 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.260 1.700 ;
        RECT  2.240 0.785 5.300 1.125 ;
        RECT  4.280 1.360 5.365 1.700 ;
        RECT  5.135 1.930 5.620 2.270 ;
        RECT  5.135 1.360 5.365 3.140 ;
        RECT  2.025 3.470 5.145 3.700 ;
        RECT  2.025 2.860 2.365 3.910 ;
        RECT  4.805 2.910 5.145 3.910 ;
        RECT  5.595 1.360 6.080 1.700 ;
        RECT  5.850 1.945 6.790 2.285 ;
        RECT  5.850 1.360 6.080 3.545 ;
        RECT  5.540 3.315 5.880 4.180 ;
        RECT  0.860 1.360 2.50 1.700 ;
        RECT  2.240 0.785 4.60 1.125 ;
        RECT  2.025 3.470 4.80 3.700 ;
    END
END ON222X4

MACRO ON222X2
    CLASS CORE ;
    FOREIGN ON222X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 3.430 3.675 4.025 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 3.430 4.325 4.030 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.435 2.120 4.935 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.150 3.430 5.545 4.040 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.080 6.210 2.630 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.685 2.640 1.135 3.560 ;
        RECT  0.685 1.250 1.080 1.590 ;
        RECT  0.685 1.250 0.915 3.560 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.800 3.430 7.435 3.895 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.775 3.430 6.115 5.280 ;
        RECT  2.790 2.740 3.130 3.080 ;
        RECT  2.790 2.740 3.075 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  3.590 -0.400 3.950 1.045 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.150 2.070 2.400 2.410 ;
        RECT  2.060 1.250 2.400 3.560 ;
        RECT  2.830 1.360 3.170 1.800 ;
        RECT  2.830 1.460 5.810 1.800 ;
        RECT  6.280 1.280 6.755 1.620 ;
        RECT  2.630 2.070 3.745 2.410 ;
        RECT  3.515 2.070 3.745 3.200 ;
        RECT  6.475 1.280 6.755 3.200 ;
        RECT  3.515 2.860 7.380 3.200 ;
        RECT  4.910 0.710 7.380 1.050 ;
        RECT  2.830 1.460 4.50 1.800 ;
        RECT  3.515 2.860 6.70 3.200 ;
        RECT  4.910 0.710 6.70 1.050 ;
    END
END ON222X2

MACRO ON222X1
    CLASS CORE ;
    FOREIGN ON222X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.345 2.120 1.765 3.240 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.795 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.285 3.240 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 4.915 2.680 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.394  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.815 3.470 5.545 3.910 ;
        RECT  4.815 2.910 5.495 3.910 ;
        RECT  5.215 1.360 5.495 3.910 ;
        RECT  4.305 1.360 5.495 1.700 ;
        RECT  2.025 3.530 5.545 3.760 ;
        RECT  2.025 2.860 2.365 3.760 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.965 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.535 3.990 3.875 5.280 ;
        RECT  0.380 2.860 0.720 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  1.550 -0.400 1.890 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.865 1.360 3.275 1.700 ;
        RECT  2.250 0.800 5.330 1.130 ;
        RECT  0.865 1.360 2.30 1.700 ;
        RECT  2.250 0.800 4.20 1.130 ;
    END
END ON222X1

MACRO ON222X0
    CLASS CORE ;
    FOREIGN ON222X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.435 4.285 3.240 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.480 0.505 3.240 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.900 1.135 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.305 2.785 1.845 3.240 ;
        RECT  1.410 2.760 1.750 3.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.500 0.630 2.910 0.860 ;
        RECT  2.160 2.250 2.445 2.820 ;
        RECT  2.015 2.250 2.445 2.630 ;
        RECT  1.500 2.250 2.445 2.505 ;
        RECT  1.500 0.630 1.730 2.505 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.135 2.010 3.655 2.630 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.156  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 3.470 3.880 3.850 ;
        RECT  2.675 1.550 3.190 1.780 ;
        RECT  2.675 1.550 2.905 3.850 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  2.440 4.170 2.780 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  0.645 -0.400 0.985 1.475 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.050 1.090 3.995 1.320 ;
        RECT  3.650 1.035 3.995 1.375 ;
        RECT  2.050 1.090 2.390 1.470 ;
    END
END ON222X0

MACRO ON221X4
    CLASS CORE ;
    FOREIGN ON221X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.340 2.120 1.765 3.240 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.780 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.160 2.120 3.675 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.366  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.080 4.275 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.960 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 0.780 8.065 3.960 ;
        RECT  6.390 2.050 8.065 2.280 ;
        RECT  6.230 2.640 6.620 3.750 ;
        RECT  6.390 1.110 6.620 3.750 ;
        RECT  6.230 1.110 6.620 1.450 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.950 2.640 7.290 5.280 ;
        RECT  5.670 4.160 6.010 5.280 ;
        RECT  3.410 3.430 3.750 5.280 ;
        RECT  0.375 2.860 0.715 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.950 -0.400 7.290 1.700 ;
        RECT  5.680 -0.400 6.020 0.710 ;
        RECT  1.540 -0.400 1.880 1.125 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.860 1.360 3.260 1.700 ;
        RECT  2.240 0.785 3.940 1.125 ;
        RECT  4.320 0.785 4.735 1.125 ;
        RECT  4.505 1.930 4.990 2.270 ;
        RECT  4.505 0.785 4.735 3.200 ;
        RECT  2.025 2.860 4.735 3.200 ;
        RECT  2.025 2.860 2.365 3.910 ;
        RECT  4.965 1.360 5.450 1.700 ;
        RECT  5.220 1.945 6.160 2.285 ;
        RECT  5.220 1.360 5.450 3.585 ;
        RECT  4.910 3.355 5.250 4.180 ;
        RECT  0.860 1.360 2.60 1.700 ;
        RECT  2.025 2.860 3.80 3.200 ;
    END
END ON221X4

MACRO ON221X2
    CLASS CORE ;
    FOREIGN ON221X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 3.430 3.675 4.090 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 3.430 4.325 4.030 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.435 2.120 4.935 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 3.430 5.545 4.045 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.685 2.640 1.135 3.560 ;
        RECT  0.685 1.250 1.080 1.590 ;
        RECT  0.685 1.250 0.920 3.560 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.770 2.095 6.230 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.775 3.560 6.115 5.280 ;
        RECT  2.790 2.740 3.130 3.080 ;
        RECT  2.790 2.740 3.075 5.280 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  3.520 -0.400 3.880 1.045 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.060 1.250 2.400 1.590 ;
        RECT  1.150 2.070 2.290 2.410 ;
        RECT  2.060 1.250 2.290 3.560 ;
        RECT  2.060 2.640 2.400 3.560 ;
        RECT  2.760 1.360 3.100 1.800 ;
        RECT  2.760 1.460 4.420 1.800 ;
        RECT  5.600 1.460 5.940 1.800 ;
        RECT  2.760 1.570 5.940 1.800 ;
        RECT  4.840 0.710 5.950 1.050 ;
        RECT  4.840 0.710 5.180 1.340 ;
        RECT  6.360 0.710 6.700 1.050 ;
        RECT  2.520 2.070 3.590 2.410 ;
        RECT  3.360 2.070 3.590 3.200 ;
        RECT  6.360 2.820 6.700 3.200 ;
        RECT  6.470 0.710 6.700 3.200 ;
        RECT  3.360 2.860 6.700 3.200 ;
        RECT  2.760 1.570 4.90 1.800 ;
        RECT  3.360 2.860 5.50 3.200 ;
    END
END ON221X2

MACRO ON221X1
    CLASS CORE ;
    FOREIGN ON221X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.345 2.120 1.765 3.240 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.795 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.655 3.240 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.361  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.285 2.700 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.025 3.470 4.865 3.760 ;
        RECT  4.525 1.360 4.865 3.760 ;
        RECT  4.385 2.955 4.865 3.760 ;
        RECT  4.305 1.360 4.865 1.700 ;
        RECT  2.025 2.950 2.365 3.760 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.965 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.535 3.990 3.875 5.280 ;
        RECT  0.380 2.860 0.720 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.550 -0.400 1.890 1.130 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.865 1.360 3.275 1.700 ;
        RECT  2.250 0.800 3.960 1.130 ;
        RECT  0.865 1.360 2.60 1.700 ;
    END
END ON221X1

MACRO ON221X0
    CLASS CORE ;
    FOREIGN ON221X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.480 0.505 3.240 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 2.235 1.300 2.685 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.650 1.640 1.955 2.290 ;
        RECT  1.385 1.640 1.955 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.175  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 0.630 2.840 0.950 ;
        RECT  2.080 2.575 2.415 2.915 ;
        RECT  2.185 0.630 2.415 2.915 ;
        RECT  2.015 0.630 2.415 1.410 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.147  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.890 3.130 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.830  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.170 3.145 3.655 3.465 ;
        RECT  3.365 1.240 3.655 3.465 ;
        RECT  3.275 2.860 3.655 3.465 ;
        RECT  2.760 1.240 3.655 1.580 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.360 4.170 2.700 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  0.645 -0.400 0.985 1.475 ;
        END
    END gnd!
END ON221X0

MACRO ON21X4
    CLASS CORE ;
    FOREIGN ON21X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.100 0.670 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.329  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.095 2.395 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.100 1.765 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.331  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 0.780 6.175 3.960 ;
        RECT  4.500 2.050 6.175 2.280 ;
        RECT  4.340 2.640 4.730 3.750 ;
        RECT  4.500 1.110 4.730 3.750 ;
        RECT  4.340 1.110 4.730 1.450 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.060 2.640 5.400 5.280 ;
        RECT  3.780 4.160 4.120 5.280 ;
        RECT  2.320 3.320 2.660 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.060 -0.400 5.400 1.700 ;
        RECT  3.790 -0.400 4.130 0.710 ;
        RECT  0.900 -0.400 1.240 1.200 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.820 0.520 1.660 ;
        RECT  1.620 0.820 1.960 1.660 ;
        RECT  0.180 1.430 1.960 1.660 ;
        RECT  2.340 0.820 2.825 1.160 ;
        RECT  2.595 0.820 2.825 1.980 ;
        RECT  2.625 2.120 3.440 2.460 ;
        RECT  2.625 1.860 2.855 3.090 ;
        RECT  1.470 2.860 2.855 3.090 ;
        RECT  1.470 2.860 1.810 3.930 ;
        RECT  3.055 1.360 3.900 1.700 ;
        RECT  3.670 1.945 4.270 2.285 ;
        RECT  3.670 1.360 3.900 3.585 ;
        RECT  3.020 3.355 3.900 3.585 ;
        RECT  3.020 3.355 3.360 4.180 ;
    END
END ON21X4

MACRO ON21X2
    CLASS CORE ;
    FOREIGN ON21X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 2.250 3.705 2.760 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.640 1.240 3.560 ;
        RECT  0.755 1.250 1.240 1.590 ;
        RECT  0.755 1.250 0.985 3.560 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.490 2.250 5.130 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.875 3.460 4.350 3.980 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.790 -0.400 4.130 1.560 ;
        RECT  1.620 -0.400 1.960 1.560 ;
        RECT  0.180 -0.400 0.520 1.560 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.025 2.860 5.365 5.280 ;
        RECT  3.070 2.990 3.415 5.280 ;
        RECT  1.620 2.640 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.190 1.255 2.680 1.595 ;
        RECT  1.380 1.945 2.420 2.285 ;
        RECT  2.190 1.255 2.420 3.560 ;
        RECT  2.190 2.640 2.680 3.560 ;
        RECT  2.805 1.790 5.450 2.020 ;
        RECT  5.110 1.220 5.450 2.020 ;
        RECT  2.650 1.945 3.035 2.285 ;
        RECT  3.935 1.790 4.235 3.200 ;
        RECT  3.935 2.860 4.565 3.200 ;
        RECT  2.805 1.790 4.70 2.020 ;
    END
END ON21X2

MACRO ON21X1
    CLASS CORE ;
    FOREIGN ON21X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 2.080 1.765 3.240 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.313  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.050 2.395 2.660 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.046  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.860 3.025 3.240 ;
        RECT  1.620 3.470 2.955 3.700 ;
        RECT  2.645 1.180 2.955 3.700 ;
        RECT  2.340 1.180 2.955 1.520 ;
        RECT  1.620 3.470 1.960 3.850 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.690 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.380 3.990 2.720 5.280 ;
        RECT  0.180 3.100 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  0.900 -0.400 1.240 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.180 0.520 1.800 ;
        RECT  1.620 1.180 1.970 1.800 ;
        RECT  0.180 1.570 1.970 1.800 ;
    END
END ON21X1

MACRO ON21X0
    CLASS CORE ;
    FOREIGN ON21X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.173  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.730 0.675 3.120 ;
        RECT  0.125 2.730 0.620 3.290 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.173  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.905 3.965 1.475 4.250 ;
        RECT  0.905 3.475 1.135 4.250 ;
        RECT  0.755 3.520 1.135 3.850 ;
        RECT  0.760 3.475 1.135 3.850 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.136  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.170 1.945 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.690  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 3.315 2.405 3.655 ;
        RECT  2.175 0.710 2.405 3.655 ;
        RECT  2.000 0.710 2.405 1.490 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  1.975 4.170 2.315 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.615 -0.400 0.955 1.555 ;
        END
    END gnd!
END ON21X0

MACRO ON211X4
    CLASS CORE ;
    FOREIGN ON211X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.715 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.850 2.120 2.395 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.005 3.015 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.292  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 0.890 6.805 3.960 ;
        RECT  5.130 2.050 6.805 2.280 ;
        RECT  4.970 2.640 5.360 3.750 ;
        RECT  5.130 0.890 5.360 3.750 ;
        RECT  4.970 0.890 5.360 1.700 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.409  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.945 2.120 1.515 2.470 ;
        RECT  0.755 2.860 1.175 3.240 ;
        RECT  0.945 2.120 1.175 3.240 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 2.640 6.030 5.280 ;
        RECT  4.410 4.160 4.750 5.280 ;
        RECT  2.180 3.320 2.520 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.700 ;
        RECT  4.250 -0.400 4.590 1.240 ;
        RECT  2.770 -0.400 3.110 1.240 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.860 1.960 1.090 ;
        RECT  1.620 0.860 1.960 1.200 ;
        RECT  0.180 0.860 0.520 1.700 ;
        RECT  0.900 1.320 1.240 1.700 ;
        RECT  0.900 1.470 3.475 1.700 ;
        RECT  3.245 1.930 3.730 2.270 ;
        RECT  1.405 2.860 3.475 3.090 ;
        RECT  3.245 1.470 3.475 3.200 ;
        RECT  2.950 2.860 3.475 3.200 ;
        RECT  1.405 2.860 1.720 3.910 ;
        RECT  1.380 3.570 1.720 3.910 ;
        RECT  3.530 0.900 3.935 1.240 ;
        RECT  3.705 0.900 3.935 1.700 ;
        RECT  3.705 1.470 4.190 1.700 ;
        RECT  3.960 1.945 4.900 2.285 ;
        RECT  3.960 1.470 4.190 3.585 ;
        RECT  3.650 3.355 3.990 4.180 ;
        RECT  0.900 1.470 2.60 1.700 ;
        RECT  1.405 2.860 2.90 3.090 ;
    END
END ON211X4

MACRO ON211X2
    CLASS CORE ;
    FOREIGN ON211X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.720 3.470 4.275 3.980 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.196  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 3.430 3.030 3.980 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 2.275 5.555 2.780 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.275 4.915 2.780 ;
        RECT  4.390 2.275 4.915 2.560 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.685 2.640 1.135 3.560 ;
        RECT  0.685 1.250 1.080 1.590 ;
        RECT  0.685 1.250 0.915 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.505 3.635 4.790 5.280 ;
        RECT  3.260 2.860 3.490 5.280 ;
        RECT  2.760 2.860 3.490 3.200 ;
        RECT  1.300 3.960 1.640 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.150 -0.400 5.490 0.950 ;
        RECT  1.300 -0.400 1.640 0.720 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.060 1.250 2.400 1.590 ;
        RECT  1.150 2.070 2.290 2.410 ;
        RECT  2.060 1.250 2.290 3.560 ;
        RECT  2.060 2.640 2.400 3.560 ;
        RECT  2.760 1.300 4.455 1.585 ;
        RECT  2.760 1.300 3.100 1.700 ;
        RECT  3.320 0.630 4.915 0.950 ;
        RECT  4.685 0.630 4.915 2.045 ;
        RECT  3.910 1.815 4.915 2.045 ;
        RECT  2.520 2.070 4.140 2.410 ;
        RECT  3.910 1.815 4.140 3.240 ;
        RECT  3.910 2.835 4.250 3.240 ;
        RECT  3.910 3.010 5.380 3.240 ;
        RECT  5.150 3.010 5.380 4.250 ;
        RECT  5.150 3.930 5.490 4.250 ;
    END
END ON211X2

MACRO ON211X1
    CLASS CORE ;
    FOREIGN ON211X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.405  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 2.120 1.765 2.630 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.342  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.470 2.395 3.240 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.342  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.120 3.025 2.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.768  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 3.475 3.655 3.855 ;
        RECT  3.055 3.470 3.655 3.855 ;
        RECT  3.055 3.045 3.495 3.855 ;
        RECT  3.265 1.470 3.495 3.855 ;
        RECT  0.900 1.470 3.495 1.700 ;
        RECT  0.900 1.360 1.240 1.700 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.405  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.110 0.760 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.145 4.170 2.485 5.280 ;
        RECT  0.175 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.905 -0.400 3.255 1.240 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.880 1.960 1.110 ;
        RECT  0.180 0.880 0.520 1.220 ;
        RECT  1.620 0.880 1.960 1.220 ;
    END
END ON211X1

MACRO ON211X0
    CLASS CORE ;
    FOREIGN ON211X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.560 0.505 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.150 1.295 2.630 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.159  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 0.630 2.100 0.970 ;
        RECT  1.385 0.630 1.765 1.360 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.159  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.460 2.785 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.924  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.095 3.025 3.850 ;
        RECT  1.170 3.095 3.025 3.435 ;
        RECT  1.525 1.590 1.755 3.435 ;
        RECT  0.635 1.590 1.755 1.820 ;
        RECT  0.635 1.130 0.975 1.820 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.970 4.170 2.310 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 1.700 ;
        END
    END gnd!
END ON211X0

MACRO OA33X4
    CLASS CORE ;
    FOREIGN OA33X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.070 3.030 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 2.060 3.675 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.020 4.305 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 5.070 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.485 2.860 6.175 3.240 ;
        RECT  5.485 2.120 5.825 3.240 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.170 2.120 6.805 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.298  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.470 3.550 1.960 3.890 ;
        RECT  1.470 2.640 1.905 3.890 ;
        RECT  1.470 1.110 1.905 1.450 ;
        RECT  1.470 1.110 1.700 3.890 ;
        RECT  0.125 2.160 1.700 2.410 ;
        RECT  0.125 0.795 0.520 3.890 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 2.860 6.750 5.280 ;
        RECT  2.340 3.320 2.680 5.280 ;
        RECT  0.900 2.640 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  3.620 -0.400 3.960 0.665 ;
        RECT  2.180 -0.400 2.520 0.665 ;
        RECT  0.900 -0.400 1.240 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.900 1.360 6.060 1.700 ;
        RECT  5.030 0.785 6.750 1.125 ;
        RECT  2.135 0.895 6.750 1.125 ;
        RECT  1.930 2.070 2.365 2.410 ;
        RECT  2.135 0.895 2.365 3.090 ;
        RECT  2.135 2.860 4.710 3.090 ;
        RECT  4.370 2.860 4.710 4.160 ;
        RECT  2.900 1.360 5.70 1.700 ;
        RECT  2.135 0.895 5.60 1.125 ;
        RECT  2.135 2.860 3.70 3.090 ;
    END
END OA33X4

MACRO OA33X2
    CLASS CORE ;
    FOREIGN OA33X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 3.445 2.400 4.085 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.120 3.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.190 3.470 3.655 4.080 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.805 2.120 4.305 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 3.460 4.925 4.085 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.115 2.085 5.620 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.640 1.150 3.565 ;
        RECT  0.750 1.240 1.150 1.580 ;
        RECT  0.750 1.240 1.060 3.565 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.590 3.430 5.930 5.280 ;
        RECT  1.530 2.855 1.870 3.195 ;
        RECT  1.530 2.855 1.785 5.280 ;
        RECT  0.250 4.020 0.590 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.570 -0.400 3.120 0.880 ;
        RECT  0.250 -0.400 0.590 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.220 1.320 3.880 1.660 ;
        RECT  5.060 1.320 5.400 1.660 ;
        RECT  2.220 1.430 5.400 1.660 ;
        RECT  4.300 0.860 6.120 1.090 ;
        RECT  4.300 0.860 4.645 1.200 ;
        RECT  5.780 0.860 6.120 1.700 ;
        RECT  1.290 1.890 2.335 2.230 ;
        RECT  2.100 1.890 2.335 3.200 ;
        RECT  5.890 0.860 6.120 3.200 ;
        RECT  2.100 2.860 6.120 3.200 ;
        RECT  2.220 1.430 4.60 1.660 ;
        RECT  2.100 2.860 5.80 3.200 ;
    END
END OA33X2

MACRO OA33X1
    CLASS CORE ;
    FOREIGN OA33X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.090 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.110 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 3.465 4.290 4.105 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.485 2.085 4.935 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.555 ;
        RECT  0.120 1.265 0.520 1.700 ;
        RECT  0.120 1.265 0.410 3.555 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.960 3.470 5.300 5.280 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  0.900 2.860 1.155 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.550 1.360 4.610 1.700 ;
        RECT  3.670 0.630 5.395 0.950 ;
        RECT  5.055 0.630 5.395 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  5.165 0.630 5.395 3.200 ;
        RECT  1.470 2.860 5.395 3.200 ;
        RECT  1.550 1.360 3.30 1.700 ;
        RECT  1.470 2.860 4.40 3.200 ;
    END
END OA33X1

MACRO OA33X0
    CLASS CORE ;
    FOREIGN OA33X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.995 2.395 2.630 ;
        RECT  1.695 1.995 2.395 2.335 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.370 3.470 3.025 3.855 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.950 2.185 3.655 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.640 3.470 4.340 3.840 ;
        RECT  3.640 3.470 3.980 3.985 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.510 2.355 4.915 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.510 ;
        RECT  0.125 2.760 0.520 3.090 ;
        RECT  0.125 1.030 0.520 1.510 ;
        RECT  0.125 1.030 0.455 3.090 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.330 3.470 1.850 3.975 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.215 4.070 4.555 5.280 ;
        RECT  0.725 3.940 1.065 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  0.245 -0.400 1.075 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.620 1.355 4.260 1.665 ;
        RECT  2.620 0.885 2.960 1.765 ;
        RECT  1.315 1.425 2.960 1.765 ;
        RECT  3.320 0.630 4.860 0.970 ;
        RECT  4.630 0.630 4.860 2.125 ;
        RECT  3.970 1.895 4.860 2.125 ;
        RECT  3.970 1.895 4.200 3.215 ;
        RECT  0.825 2.875 4.200 3.215 ;
        RECT  0.825 2.875 1.055 3.710 ;
        RECT  0.460 3.410 1.055 3.710 ;
        RECT  0.825 2.875 3.60 3.215 ;
    END
END OA33X0

MACRO OA333X1
    CLASS CORE ;
    FOREIGN OA333X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.120 6.940 2.630 ;
        END
    END J
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.090 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 3.465 4.290 4.090 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.485 2.085 4.935 2.630 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.085 5.580 2.630 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.860 ;
        RECT  0.120 1.265 0.520 1.605 ;
        RECT  0.120 1.265 0.410 3.860 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 3.470 6.260 3.995 ;
        END
    END H
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.090 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  4.960 3.470 5.300 5.280 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  0.900 2.860 1.155 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.550 1.360 4.610 1.700 ;
        RECT  3.670 0.630 6.620 0.950 ;
        RECT  5.670 1.360 7.420 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  7.170 1.360 7.420 3.200 ;
        RECT  1.470 2.860 7.420 3.200 ;
        RECT  1.550 1.360 3.70 1.700 ;
        RECT  3.670 0.630 5.60 0.950 ;
        RECT  1.470 2.860 6.60 3.200 ;
    END
END OA333X1

MACRO OA333X0
    CLASS CORE ;
    FOREIGN OA333X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.700 1.995 2.395 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.370 3.470 3.025 4.010 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.100 3.655 2.635 ;
        RECT  2.970 2.100 3.655 2.525 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.640 3.470 4.285 3.850 ;
        RECT  3.640 3.470 3.980 4.010 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.260 2.170 4.915 2.630 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.970 3.470 5.545 4.010 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.630 0.520 3.125 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.605 1.865 6.175 2.630 ;
        END
    END H
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.035 3.470 6.805 3.865 ;
        END
    END J
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 3.470 1.830 4.010 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  0.980 -0.400 2.320 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.215 4.080 4.555 5.280 ;
        RECT  0.780 3.900 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.680 0.885 3.020 1.765 ;
        RECT  1.380 1.425 4.320 1.765 ;
        RECT  3.380 0.665 6.350 1.005 ;
        RECT  6.010 0.665 6.350 1.470 ;
        RECT  5.145 1.300 5.550 1.635 ;
        RECT  5.145 1.300 5.375 3.240 ;
        RECT  0.830 2.900 6.655 3.240 ;
        RECT  0.830 2.900 1.060 3.670 ;
        RECT  0.460 3.355 1.060 3.670 ;
        RECT  1.380 1.425 3.90 1.765 ;
        RECT  3.380 0.665 5.70 1.005 ;
        RECT  0.830 2.900 5.00 3.240 ;
    END
END OA333X0

MACRO OA332X1
    CLASS CORE ;
    FOREIGN OA332X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.090 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 3.465 4.290 4.105 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.485 2.085 4.935 2.630 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.080 5.580 2.630 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.860 ;
        RECT  0.120 1.265 0.520 1.605 ;
        RECT  0.120 1.265 0.410 3.860 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.090 ;
        END
    END A
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 3.470 6.260 3.995 ;
        END
    END H
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.960 3.470 5.300 5.280 ;
        RECT  0.900 2.865 1.240 3.205 ;
        RECT  0.900 2.865 1.155 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.550 1.360 4.610 1.700 ;
        RECT  3.670 0.630 6.620 0.950 ;
        RECT  5.670 1.360 6.745 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  6.485 1.360 6.745 3.200 ;
        RECT  1.470 2.860 6.745 3.200 ;
        RECT  1.550 1.360 3.30 1.700 ;
        RECT  3.670 0.630 5.20 0.950 ;
        RECT  1.470 2.860 5.70 3.200 ;
    END
END OA332X1

MACRO OA332X0
    CLASS CORE ;
    FOREIGN OA332X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.965 2.395 2.630 ;
        RECT  1.650 1.965 2.395 2.285 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.370 3.670 3.025 4.010 ;
        RECT  2.645 3.380 3.025 4.010 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.100 3.655 2.635 ;
        RECT  2.955 2.100 3.655 2.525 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.640 3.460 4.285 3.850 ;
        RECT  3.640 3.460 3.980 4.010 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.260 2.150 4.880 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.408  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.030 0.785 1.510 ;
        RECT  0.125 1.030 0.520 3.150 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.570 2.250 6.175 2.630 ;
        RECT  5.570 1.945 5.860 2.630 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.760 3.470 5.545 3.865 ;
        END
    END G
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.380 1.785 3.960 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  0.445 -0.400 2.320 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.215 4.080 4.555 5.280 ;
        RECT  0.780 3.950 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.545 0.885 2.885 1.710 ;
        RECT  1.245 1.425 4.185 1.710 ;
        RECT  1.245 1.425 1.570 1.745 ;
        RECT  3.845 1.425 4.185 1.815 ;
        RECT  3.245 0.840 4.785 1.180 ;
        RECT  5.110 1.210 5.585 1.550 ;
        RECT  5.110 1.210 5.340 3.150 ;
        RECT  2.650 2.810 2.990 3.150 ;
        RECT  5.110 2.860 6.025 3.150 ;
        RECT  0.925 2.865 6.025 3.150 ;
        RECT  0.925 2.865 1.155 3.720 ;
        RECT  0.460 3.380 1.155 3.720 ;
        RECT  1.245 1.425 3.70 1.710 ;
        RECT  0.925 2.865 5.60 3.150 ;
    END
END OA332X0

MACRO OA331X1
    CLASS CORE ;
    FOREIGN OA331X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.090 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.860 ;
        RECT  0.120 1.265 0.520 1.605 ;
        RECT  0.120 1.265 0.410 3.860 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.995 5.580 2.630 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.485 2.085 4.935 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 3.465 4.290 4.090 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.960 3.470 5.300 5.280 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  0.900 2.860 1.155 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.550 1.360 4.610 1.700 ;
        RECT  3.670 0.630 5.290 0.950 ;
        RECT  5.670 1.360 6.125 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  5.845 1.360 6.125 3.200 ;
        RECT  1.470 2.860 6.125 3.200 ;
        RECT  1.550 1.360 3.50 1.700 ;
        RECT  1.470 2.860 5.80 3.200 ;
    END
END OA331X1

MACRO OA331X0
    CLASS CORE ;
    FOREIGN OA331X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.695 1.995 2.395 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.370 3.470 3.025 3.850 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.100 3.655 2.630 ;
        RECT  2.950 2.100 3.655 2.525 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.640 3.470 4.285 3.850 ;
        RECT  3.640 3.470 3.980 3.960 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.135 2.095 4.915 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.408  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.510 ;
        RECT  0.125 2.760 0.520 3.075 ;
        RECT  0.125 1.030 0.520 1.510 ;
        RECT  0.125 1.030 0.455 3.075 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.735 3.470 5.545 3.850 ;
        END
    END G
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.350 3.470 1.915 3.865 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  0.435 -0.400 2.185 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.215 4.080 4.555 5.280 ;
        RECT  0.780 3.840 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.545 0.885 2.885 1.765 ;
        RECT  1.245 1.425 4.185 1.765 ;
        RECT  3.245 0.710 4.785 1.050 ;
        RECT  5.145 0.710 5.490 3.190 ;
        RECT  0.825 2.860 5.490 3.190 ;
        RECT  0.825 2.860 1.055 3.610 ;
        RECT  0.460 3.305 1.055 3.610 ;
        RECT  1.245 1.425 3.20 1.765 ;
        RECT  0.825 2.860 4.30 3.190 ;
    END
END OA331X0

MACRO OA32X4
    CLASS CORE ;
    FOREIGN OA32X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.070 3.030 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 2.060 3.675 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.020 4.305 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.471  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.120 5.070 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.485 2.120 6.175 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.298  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.470 3.550 1.960 3.890 ;
        RECT  1.470 2.640 1.905 3.890 ;
        RECT  1.470 1.110 1.905 1.450 ;
        RECT  1.470 1.110 1.700 3.890 ;
        RECT  0.125 2.160 1.700 2.410 ;
        RECT  0.125 0.795 0.520 3.890 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.720 2.860 6.060 5.280 ;
        RECT  2.340 3.320 2.680 5.280 ;
        RECT  0.900 2.640 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  3.620 -0.400 3.960 0.665 ;
        RECT  2.180 -0.400 2.520 0.665 ;
        RECT  0.900 -0.400 1.240 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  5.030 0.785 5.375 1.125 ;
        RECT  2.135 0.895 5.375 1.125 ;
        RECT  1.930 2.070 2.365 2.410 ;
        RECT  2.135 0.895 2.365 3.090 ;
        RECT  2.135 2.860 4.710 3.090 ;
        RECT  4.370 2.860 4.710 4.160 ;
        RECT  2.900 1.360 6.060 1.700 ;
        RECT  2.135 0.895 4.20 1.125 ;
        RECT  2.135 2.860 3.50 3.090 ;
        RECT  2.900 1.360 5.10 1.700 ;
    END
END OA32X4

MACRO OA32X2
    CLASS CORE ;
    FOREIGN OA32X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 3.445 2.400 4.085 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.120 3.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.190 3.470 3.655 4.080 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 3.460 4.920 4.085 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.805 2.120 4.305 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.640 1.150 3.570 ;
        RECT  0.750 1.240 1.150 1.580 ;
        RECT  0.750 1.240 1.060 3.570 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 2.640 5.490 5.280 ;
        RECT  1.530 2.920 1.870 3.260 ;
        RECT  1.530 2.920 1.785 5.280 ;
        RECT  0.250 4.020 0.590 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  1.570 -0.400 3.120 0.880 ;
        RECT  0.250 -0.400 0.590 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  4.300 1.320 4.765 1.660 ;
        RECT  1.290 1.890 2.335 2.230 ;
        RECT  2.100 1.890 2.335 3.200 ;
        RECT  4.535 1.320 4.765 3.200 ;
        RECT  2.100 2.860 4.765 3.200 ;
        RECT  3.540 0.860 5.400 1.090 ;
        RECT  3.540 0.860 3.880 1.660 ;
        RECT  2.220 1.320 3.880 1.660 ;
        RECT  5.060 0.860 5.400 1.660 ;
        RECT  2.100 2.860 3.40 3.200 ;
    END
END OA32X2

MACRO OA32X1
    CLASS CORE ;
    FOREIGN OA32X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.085 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.535 ;
        RECT  0.120 1.265 0.520 1.700 ;
        RECT  0.120 1.265 0.410 3.535 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 3.465 4.285 4.085 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.085 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.515 2.660 4.855 5.280 ;
        RECT  0.900 2.865 1.240 3.205 ;
        RECT  0.900 2.865 1.155 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.630 1.360 4.145 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  3.915 1.360 4.145 3.200 ;
        RECT  1.470 2.860 4.145 3.200 ;
        RECT  2.910 0.900 4.730 1.130 ;
        RECT  4.375 0.900 4.730 1.690 ;
        RECT  2.910 0.900 3.250 1.700 ;
        RECT  1.550 1.360 3.250 1.700 ;
        RECT  1.470 2.860 3.80 3.200 ;
    END
END OA32X1

MACRO OA32X0
    CLASS CORE ;
    FOREIGN OA32X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.650 3.470 1.990 4.070 ;
        RECT  1.385 3.470 1.990 3.850 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.945 2.610 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.440 3.220 3.850 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.060 3.835 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.460 ;
        RECT  0.125 2.870 0.520 3.185 ;
        RECT  0.125 1.030 0.520 1.460 ;
        RECT  0.125 1.030 0.455 3.185 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.725 2.250 1.135 2.630 ;
        RECT  0.725 1.690 1.015 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.630 3.655 3.970 5.280 ;
        RECT  0.780 4.040 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  0.445 -0.400 2.185 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.655 0.885 2.995 1.710 ;
        RECT  1.315 1.425 2.995 1.710 ;
        RECT  1.315 1.425 1.655 1.765 ;
        RECT  3.355 1.255 4.295 1.595 ;
        RECT  4.065 1.255 4.295 3.210 ;
        RECT  0.750 2.870 4.295 3.210 ;
        RECT  0.750 2.870 0.980 3.810 ;
        RECT  0.460 3.505 0.980 3.810 ;
        RECT  0.750 2.870 3.40 3.210 ;
    END
END OA32X0

MACRO OA322X1
    CLASS CORE ;
    FOREIGN OA322X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 3.470 6.260 3.995 ;
        END
    END G
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.090 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.860 ;
        RECT  0.120 1.245 0.520 1.585 ;
        RECT  0.120 1.245 0.350 3.860 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.995 5.580 2.630 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 3.465 4.285 4.105 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.175 2.120 3.675 2.630 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.165 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.515 3.470 5.300 5.280 ;
        RECT  0.900 2.920 1.240 3.260 ;
        RECT  0.900 2.920 1.155 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.550 1.360 1.890 1.700 ;
        RECT  2.910 1.360 3.250 1.700 ;
        RECT  4.270 1.360 4.610 1.700 ;
        RECT  1.550 1.470 4.610 1.700 ;
        RECT  3.670 0.630 6.580 0.950 ;
        RECT  5.630 1.360 6.040 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  5.810 1.360 6.040 3.200 ;
        RECT  1.470 2.860 6.625 3.200 ;
        RECT  1.550 1.470 3.40 1.700 ;
        RECT  3.670 0.630 5.30 0.950 ;
        RECT  1.470 2.860 5.20 3.200 ;
    END
END OA322X1

MACRO OA322X0
    CLASS CORE ;
    FOREIGN OA322X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.695 1.960 2.395 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.370 3.470 3.025 3.865 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.930 2.095 3.655 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.600 3.420 4.285 3.850 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.408  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.510 ;
        RECT  0.125 2.760 0.520 3.075 ;
        RECT  0.125 1.030 0.520 1.510 ;
        RECT  0.125 1.030 0.455 3.075 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.870 3.470 5.545 3.865 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.200 2.030 4.915 2.630 ;
        END
    END F
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 3.420 1.815 3.955 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  0.445 -0.400 2.185 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.920 4.080 4.260 5.280 ;
        RECT  0.780 3.840 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.545 0.885 2.885 1.710 ;
        RECT  1.245 1.425 2.885 1.710 ;
        RECT  1.245 1.425 1.570 1.750 ;
        RECT  3.245 0.715 4.385 1.055 ;
        RECT  3.245 0.715 3.585 1.765 ;
        RECT  4.735 1.210 5.490 1.550 ;
        RECT  5.215 1.210 5.490 3.190 ;
        RECT  0.830 2.860 5.490 3.190 ;
        RECT  0.830 2.860 1.060 3.610 ;
        RECT  0.460 3.305 1.060 3.610 ;
        RECT  0.830 2.860 4.50 3.190 ;
    END
END OA322X0

MACRO OA321X4
    CLASS CORE ;
    FOREIGN OA321X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.080 3.755 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.260 2.080 4.915 2.630 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.080 7.510 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 2.020 5.545 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.055 6.200 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.254  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.615 3.550 1.960 3.890 ;
        RECT  1.615 1.130 1.960 1.470 ;
        RECT  1.615 2.665 1.955 3.890 ;
        RECT  1.615 1.130 1.845 3.890 ;
        RECT  0.125 1.985 1.845 2.235 ;
        RECT  0.125 1.130 0.520 3.890 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.020 3.045 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.910 3.320 7.250 5.280 ;
        RECT  6.050 3.320 6.390 5.280 ;
        RECT  2.425 3.320 2.765 5.280 ;
        RECT  0.900 2.640 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  3.780 -0.400 4.120 1.300 ;
        RECT  2.340 -0.400 2.680 1.470 ;
        RECT  0.900 -0.400 1.240 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.060 1.160 3.400 1.760 ;
        RECT  4.555 1.160 4.895 1.760 ;
        RECT  6.050 1.360 6.390 1.760 ;
        RECT  3.060 1.530 6.390 1.760 ;
        RECT  5.330 0.900 7.110 1.130 ;
        RECT  5.330 0.900 5.670 1.300 ;
        RECT  6.770 0.900 7.110 1.500 ;
        RECT  7.490 1.160 7.970 1.500 ;
        RECT  2.075 2.120 2.415 2.460 ;
        RECT  2.185 2.120 2.415 3.090 ;
        RECT  2.185 2.860 7.970 3.090 ;
        RECT  4.555 2.860 4.895 4.160 ;
        RECT  7.740 1.160 7.970 4.160 ;
        RECT  7.630 2.860 7.970 4.160 ;
        RECT  3.060 1.530 5.00 1.760 ;
        RECT  2.185 2.860 6.40 3.090 ;
    END
END OA321X4

MACRO OA321X2
    CLASS CORE ;
    FOREIGN OA321X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.540 2.190 3.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.190 3.470 3.655 4.250 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.740 2.190 4.340 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 3.465 4.915 4.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.710 2.840 1.135 3.760 ;
        RECT  0.710 1.240 1.080 1.580 ;
        RECT  0.710 1.240 0.940 3.760 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 3.450 2.395 4.250 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.160 2.080 5.605 2.630 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.145 4.160 5.480 5.280 ;
        RECT  1.460 2.840 1.785 3.180 ;
        RECT  1.460 2.840 1.780 5.280 ;
        RECT  0.180 4.160 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.500 -0.400 2.960 0.880 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.060 1.320 5.040 1.660 ;
        RECT  4.700 1.320 5.040 1.820 ;
        RECT  4.140 0.640 5.780 0.990 ;
        RECT  4.140 0.640 4.480 1.080 ;
        RECT  5.440 1.360 6.080 1.700 ;
        RECT  1.170 2.265 2.245 2.605 ;
        RECT  2.015 2.265 2.245 3.200 ;
        RECT  2.015 2.860 6.080 3.200 ;
        RECT  5.850 1.360 6.080 3.760 ;
        RECT  5.740 2.860 6.080 3.760 ;
        RECT  2.060 1.320 4.80 1.660 ;
        RECT  2.015 2.860 5.40 3.200 ;
    END
END OA321X2

MACRO OA321X1
    CLASS CORE ;
    FOREIGN OA321X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.470 1.780 4.085 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.700 0.520 3.620 ;
        RECT  0.125 1.265 0.520 1.605 ;
        RECT  0.125 1.265 0.360 3.620 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.910 3.470 5.545 3.940 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.180 4.400 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.155 2.165 3.670 2.630 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.470 3.060 4.070 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.975 2.175 2.510 2.630 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  0.940 -0.400 2.400 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.285 3.460 4.625 5.280 ;
        RECT  0.900 2.920 1.240 3.260 ;
        RECT  0.900 2.920 1.155 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.500 1.360 4.480 1.700 ;
        RECT  4.140 1.360 4.480 1.750 ;
        RECT  3.580 0.670 4.770 1.040 ;
        RECT  0.590 1.940 1.700 2.280 ;
        RECT  1.470 1.940 1.700 3.230 ;
        RECT  5.150 0.710 5.490 3.230 ;
        RECT  1.470 2.890 5.490 3.230 ;
        RECT  1.500 1.360 3.90 1.700 ;
        RECT  1.470 2.890 4.40 3.230 ;
    END
END OA321X1

MACRO OA321X0
    CLASS CORE ;
    FOREIGN OA321X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.650 3.470 1.990 3.960 ;
        RECT  1.385 3.470 1.990 3.850 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.000 2.635 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.470 3.220 3.910 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.045 3.890 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.030 0.785 1.370 ;
        RECT  0.125 2.760 0.520 3.075 ;
        RECT  0.125 1.030 0.455 3.075 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.240 3.470 4.915 3.865 ;
        END
    END F
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.725 2.250 1.135 2.630 ;
        RECT  0.725 1.690 1.015 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.670 3.540 4.010 5.280 ;
        RECT  0.780 3.930 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.110 -0.400 2.185 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.655 0.885 2.995 1.765 ;
        RECT  1.245 1.425 4.295 1.765 ;
        RECT  4.345 0.630 4.860 0.965 ;
        RECT  4.525 0.630 4.860 3.190 ;
        RECT  0.840 2.860 4.860 3.190 ;
        RECT  0.840 2.860 1.070 3.700 ;
        RECT  0.460 3.395 1.070 3.700 ;
        RECT  1.245 1.425 3.90 1.765 ;
        RECT  0.840 2.860 3.30 3.190 ;
    END
END OA321X0

MACRO OA31X4
    CLASS CORE ;
    FOREIGN OA31X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.020 3.045 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.020 3.675 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.060 4.305 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.110 5.005 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.332  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.515 3.550 1.960 3.890 ;
        RECT  1.515 1.110 1.960 1.450 ;
        RECT  1.515 2.640 1.955 3.890 ;
        RECT  1.515 1.110 1.745 3.890 ;
        RECT  0.125 2.160 1.745 2.410 ;
        RECT  0.125 0.795 0.520 3.890 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.135 3.320 5.475 5.280 ;
        RECT  2.405 3.320 2.745 5.280 ;
        RECT  0.900 2.640 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.660 -0.400 4.000 1.300 ;
        RECT  2.180 -0.400 2.520 0.710 ;
        RECT  0.900 -0.400 1.240 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.940 1.160 3.280 1.760 ;
        RECT  4.380 1.160 4.720 1.760 ;
        RECT  2.940 1.530 4.720 1.760 ;
        RECT  5.135 1.160 5.480 1.500 ;
        RECT  1.975 2.070 2.415 2.410 ;
        RECT  2.185 2.070 2.415 3.090 ;
        RECT  5.250 1.160 5.480 3.090 ;
        RECT  2.185 2.860 5.480 3.090 ;
        RECT  4.320 2.860 4.660 4.160 ;
        RECT  2.185 2.860 4.20 3.090 ;
    END
END OA31X4

MACRO OA31X2
    CLASS CORE ;
    FOREIGN OA31X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 3.445 2.400 4.085 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.120 3.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.190 3.470 3.655 4.080 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 3.460 4.290 4.085 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.640 1.150 3.560 ;
        RECT  0.750 1.240 1.150 1.580 ;
        RECT  0.750 1.240 1.060 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.520 2.640 4.860 5.280 ;
        RECT  1.530 2.920 1.870 3.260 ;
        RECT  1.530 2.920 1.785 5.280 ;
        RECT  0.250 4.020 0.590 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.570 -0.400 3.120 0.880 ;
        RECT  0.250 -0.400 0.590 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.220 1.320 3.880 1.660 ;
        RECT  1.290 1.890 2.400 2.230 ;
        RECT  4.295 1.320 4.635 2.300 ;
        RECT  3.685 2.070 4.635 2.300 ;
        RECT  2.165 1.890 2.400 3.200 ;
        RECT  3.685 2.070 3.915 3.200 ;
        RECT  2.165 2.860 3.915 3.200 ;
    END
END OA31X2

MACRO OA31X1
    CLASS CORE ;
    FOREIGN OA31X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.120 2.505 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 3.470 3.025 4.035 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 3.470 3.655 4.035 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.640 0.520 3.550 ;
        RECT  0.120 1.265 0.520 1.700 ;
        RECT  0.120 1.265 0.410 3.550 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.450 1.765 4.035 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.885 2.640 4.225 5.280 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  0.900 2.860 1.155 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  0.940 -0.400 2.490 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.550 1.360 3.250 1.700 ;
        RECT  0.640 1.940 1.770 2.280 ;
        RECT  3.630 1.360 3.970 2.330 ;
        RECT  2.985 1.990 3.970 2.330 ;
        RECT  1.470 1.940 1.770 3.200 ;
        RECT  2.985 1.990 3.305 3.200 ;
        RECT  1.470 2.860 3.305 3.200 ;
    END
END OA31X1

MACRO OA31X0
    CLASS CORE ;
    FOREIGN OA31X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 3.470 1.885 3.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.140 2.535 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.555 3.430 3.095 3.845 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.516  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.460 ;
        RECT  0.125 2.750 0.520 3.065 ;
        RECT  0.125 1.030 0.520 1.460 ;
        RECT  0.125 1.030 0.485 3.065 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.725 2.250 1.135 2.630 ;
        RECT  0.725 1.690 1.015 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.075 4.075 3.415 5.280 ;
        RECT  0.780 3.920 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  1.055 -0.400 2.335 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.645 1.315 2.985 1.765 ;
        RECT  1.245 1.425 2.985 1.765 ;
        RECT  1.245 1.425 1.590 1.835 ;
        RECT  3.245 0.630 3.585 0.970 ;
        RECT  3.345 0.630 3.585 3.180 ;
        RECT  0.815 2.860 3.585 3.180 ;
        RECT  0.815 2.860 1.045 3.690 ;
        RECT  0.460 3.385 1.045 3.690 ;
        RECT  0.815 2.860 2.80 3.180 ;
    END
END OA31X0

MACRO OA311X4
    CLASS CORE ;
    FOREIGN OA311X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.020 3.675 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.020 4.305 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.770 2.045 6.185 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.080 5.080 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.254  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.515 3.550 1.960 3.890 ;
        RECT  1.515 1.130 1.960 1.470 ;
        RECT  1.515 2.690 1.955 3.890 ;
        RECT  1.515 1.130 1.745 3.890 ;
        RECT  0.125 1.985 1.745 2.235 ;
        RECT  0.125 1.130 0.520 3.890 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.020 3.045 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.020 3.320 5.360 5.280 ;
        RECT  2.380 3.320 2.720 5.280 ;
        RECT  0.900 2.640 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  3.780 -0.400 4.120 1.300 ;
        RECT  2.340 -0.400 2.680 1.470 ;
        RECT  0.900 -0.400 1.240 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.060 1.160 3.400 1.760 ;
        RECT  4.500 1.160 4.840 1.760 ;
        RECT  3.060 1.530 4.840 1.760 ;
        RECT  5.310 1.160 6.080 1.500 ;
        RECT  1.975 2.120 2.415 2.460 ;
        RECT  2.185 2.120 2.415 3.090 ;
        RECT  5.310 1.160 5.540 3.090 ;
        RECT  2.185 2.860 6.125 3.090 ;
        RECT  4.300 2.860 4.640 4.160 ;
        RECT  5.740 2.860 6.125 4.160 ;
        RECT  2.185 2.860 5.60 3.090 ;
    END
END OA311X4

MACRO OA311X2
    CLASS CORE ;
    FOREIGN OA311X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.240 2.640 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 3.470 3.300 4.250 ;
        RECT  2.645 3.470 3.300 3.850 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.280 3.470 4.620 4.250 ;
        RECT  3.905 3.470 4.620 3.850 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.235 3.950 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 2.840 1.080 3.760 ;
        RECT  0.690 1.240 1.080 1.580 ;
        RECT  0.690 1.240 0.920 3.760 ;
        RECT  0.125 2.250 0.920 2.630 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.820 3.470 2.160 4.250 ;
        RECT  1.385 3.470 2.160 3.850 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.710 4.160 4.050 5.280 ;
        RECT  1.250 4.160 1.590 5.280 ;
        RECT  0.180 4.160 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.500 -0.400 2.960 0.880 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.320 0.630 3.660 1.660 ;
        RECT  2.060 1.320 3.660 1.660 ;
        RECT  4.520 1.320 4.860 1.660 ;
        RECT  1.150 2.265 1.595 2.605 ;
        RECT  1.365 2.265 1.595 3.200 ;
        RECT  4.630 1.320 4.860 3.200 ;
        RECT  1.365 2.860 4.860 3.200 ;
        RECT  1.365 2.860 3.30 3.200 ;
    END
END OA311X2

MACRO OA311X1
    CLASS CORE ;
    FOREIGN OA311X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.310 3.470 1.765 4.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.640 0.520 3.560 ;
        RECT  0.125 1.240 0.520 1.580 ;
        RECT  0.125 1.240 0.360 3.560 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.060 2.120 3.670 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 1.620 4.295 2.240 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.385 3.465 2.975 3.885 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.720 2.120 2.395 2.630 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  0.940 -0.400 2.400 0.725 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.205 3.760 3.530 5.280 ;
        RECT  0.740 3.960 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.500 1.415 3.160 1.700 ;
        RECT  3.810 0.630 4.150 1.185 ;
        RECT  0.750 0.955 4.150 1.185 ;
        RECT  0.590 2.070 0.980 2.410 ;
        RECT  0.750 0.955 0.980 3.230 ;
        RECT  0.750 2.890 4.230 3.230 ;
        RECT  3.890 2.890 4.230 4.100 ;
        RECT  0.750 0.955 3.20 1.185 ;
        RECT  0.750 2.890 3.50 3.230 ;
    END
END OA311X1

MACRO OA311X0
    CLASS CORE ;
    FOREIGN OA311X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.470 1.890 3.955 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.995 2.555 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.510 3.470 3.095 3.920 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.030 0.785 1.320 ;
        RECT  0.125 2.755 0.520 3.070 ;
        RECT  0.125 1.030 0.455 3.070 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 3.320 4.285 3.850 ;
        RECT  3.595 3.320 4.285 3.615 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.725 2.250 1.135 2.630 ;
        RECT  0.725 1.690 1.015 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.325 3.845 3.665 5.280 ;
        RECT  0.780 3.925 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.140 -0.400 2.185 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.245 1.425 2.985 1.765 ;
        RECT  3.875 1.225 4.230 3.090 ;
        RECT  0.750 2.860 4.230 3.090 ;
        RECT  0.750 2.860 2.815 3.185 ;
        RECT  0.750 2.860 0.980 3.695 ;
        RECT  0.460 3.390 0.980 3.695 ;
        RECT  0.750 2.860 3.00 3.090 ;
        RECT  0.750 2.860 1.40 3.185 ;
    END
END OA311X0

MACRO OA22X4
    CLASS CORE ;
    FOREIGN OA22X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.140 3.215 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.615 3.840 1.960 4.180 ;
        RECT  1.615 1.280 1.960 1.620 ;
        RECT  1.615 2.955 1.955 4.180 ;
        RECT  1.615 1.280 1.845 4.180 ;
        RECT  0.125 2.400 1.845 2.630 ;
        RECT  0.125 0.700 0.520 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.040 6.185 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.815 2.140 5.545 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.140 4.435 2.630 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.055 -0.400 5.395 1.240 ;
        RECT  2.195 -0.400 2.535 0.710 ;
        RECT  0.900 -0.400 1.240 1.620 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 2.860 6.120 5.280 ;
        RECT  2.340 3.320 3.480 5.280 ;
        RECT  0.900 2.930 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.445 1.280 3.955 1.620 ;
        RECT  2.075 2.410 2.415 2.750 ;
        RECT  2.185 2.410 2.415 3.090 ;
        RECT  3.445 1.280 3.675 3.090 ;
        RECT  2.185 2.860 4.795 3.090 ;
        RECT  4.455 2.860 4.795 4.180 ;
        RECT  2.895 0.820 4.675 1.050 ;
        RECT  2.895 0.820 3.235 1.160 ;
        RECT  4.335 0.820 4.675 1.700 ;
        RECT  2.895 0.820 3.215 1.700 ;
        RECT  5.780 0.820 6.120 1.700 ;
        RECT  4.335 1.470 6.120 1.700 ;
        RECT  2.185 2.860 3.60 3.090 ;
    END
END OA22X4

MACRO OA22X2
    CLASS CORE ;
    FOREIGN OA22X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.175 2.735 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.805 2.695 1.245 3.850 ;
        RECT  0.805 1.240 1.150 3.850 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.625 4.925 2.235 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.610 2.175 4.285 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.115 3.470 3.655 4.135 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.955 -0.400 4.295 1.610 ;
        RECT  1.370 -0.400 1.710 0.720 ;
        RECT  0.250 -0.400 0.590 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.520 2.805 4.860 5.280 ;
        RECT  1.625 2.860 2.500 5.280 ;
        RECT  1.625 2.845 1.930 5.280 ;
        RECT  0.180 2.695 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.385 1.270 3.345 1.610 ;
        RECT  1.385 1.270 1.725 2.220 ;
        RECT  3.115 1.270 3.345 3.240 ;
        RECT  3.115 2.900 3.700 3.240 ;
    END
END OA22X2

MACRO OA22X1
    CLASS CORE ;
    FOREIGN OA22X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 1.760 1.765 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.900 0.520 3.970 ;
        RECT  0.120 1.360 0.520 1.700 ;
        RECT  0.120 1.360 0.350 3.970 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.570 2.120 4.285 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.120 3.185 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 3.470 2.395 4.165 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.325 -0.400 3.665 1.530 ;
        RECT  0.740 -0.400 1.095 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.795 3.075 4.135 5.280 ;
        RECT  0.900 2.955 1.245 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.750 1.190 2.345 1.530 ;
        RECT  0.750 1.190 0.980 2.280 ;
        RECT  0.640 1.940 0.980 2.280 ;
        RECT  2.045 1.190 2.345 3.200 ;
        RECT  2.045 2.860 2.675 3.200 ;
    END
END OA22X1

MACRO OA22X0
    CLASS CORE ;
    FOREIGN OA22X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.050 1.320 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.455 2.070 3.930 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.955 2.645 2.295 ;
        RECT  2.015 1.640 2.395 2.295 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 0.865 3.655 1.490 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.030 0.785 1.510 ;
        RECT  0.125 2.785 0.520 3.100 ;
        RECT  0.125 1.030 0.455 3.100 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.055 3.525 3.395 5.280 ;
        RECT  0.780 3.955 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.755 -0.400 3.045 1.725 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.245 1.505 1.785 1.820 ;
        RECT  1.555 1.505 1.785 3.125 ;
        RECT  1.555 2.785 2.360 3.125 ;
        RECT  0.925 2.890 2.360 3.125 ;
        RECT  0.925 2.890 1.155 3.725 ;
        RECT  0.460 3.420 1.155 3.725 ;
    END
END OA22X0

MACRO OA222X4
    CLASS CORE ;
    FOREIGN OA222X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.580 2.100 3.045 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.880 2.055 4.305 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.055 5.565 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.990 2.095 7.445 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.055 4.935 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.440 3.320 1.960 4.160 ;
        RECT  1.440 1.290 1.840 1.630 ;
        RECT  1.440 1.290 1.670 4.160 ;
        RECT  0.180 2.250 1.670 2.630 ;
        RECT  0.180 0.700 0.520 4.160 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.120 6.300 2.630 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.720 3.320 6.060 5.280 ;
        RECT  2.340 3.320 3.355 5.280 ;
        RECT  0.900 2.910 1.210 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  3.580 -0.400 3.920 0.710 ;
        RECT  2.060 -0.400 2.400 0.710 ;
        RECT  0.940 -0.400 1.280 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.820 0.820 3.160 1.825 ;
        RECT  4.880 1.280 5.220 1.825 ;
        RECT  2.820 1.595 5.220 1.825 ;
        RECT  6.320 1.280 6.760 1.620 ;
        RECT  1.900 2.390 2.200 3.090 ;
        RECT  6.530 1.280 6.760 3.090 ;
        RECT  1.900 2.860 7.380 3.090 ;
        RECT  4.355 2.860 4.695 4.160 ;
        RECT  7.040 2.860 7.380 4.160 ;
        RECT  4.160 0.820 7.380 1.050 ;
        RECT  4.160 0.820 4.500 1.365 ;
        RECT  5.600 0.820 5.945 1.430 ;
        RECT  7.040 0.820 7.380 1.700 ;
        RECT  2.820 1.595 4.50 1.825 ;
        RECT  1.900 2.860 6.10 3.090 ;
        RECT  4.160 0.820 6.40 1.050 ;
    END
END OA222X4

MACRO OA222X2
    CLASS CORE ;
    FOREIGN OA222X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.930 2.250 2.415 2.750 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.250 3.130 2.750 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 0.900 3.675 1.440 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.765 2.250 4.285 2.720 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.250 4.935 2.750 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 3.105 1.240 4.025 ;
        RECT  0.750 0.820 1.240 1.160 ;
        RECT  0.750 0.820 1.060 4.025 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.235 5.645 2.750 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.250 3.440 4.590 5.280 ;
        RECT  1.680 3.440 2.020 5.280 ;
        RECT  0.180 3.105 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.660 -0.400 2.490 1.160 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.570 1.680 4.550 2.020 ;
        RECT  5.010 1.250 5.350 1.590 ;
        RECT  5.010 1.360 6.120 1.590 ;
        RECT  1.290 2.350 1.700 2.690 ;
        RECT  1.470 2.350 1.700 3.210 ;
        RECT  1.470 2.980 6.120 3.210 ;
        RECT  2.890 2.980 3.230 4.025 ;
        RECT  5.890 1.360 6.120 4.025 ;
        RECT  5.780 2.980 6.120 4.025 ;
        RECT  4.025 0.790 6.120 1.020 ;
        RECT  4.025 0.790 4.365 1.130 ;
        RECT  5.780 0.790 6.120 1.130 ;
        RECT  1.570 1.680 3.60 2.020 ;
        RECT  1.470 2.980 5.40 3.210 ;
        RECT  4.025 0.790 5.80 1.020 ;
    END
END OA222X2

MACRO OA222X1
    CLASS CORE ;
    FOREIGN OA222X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 3.470 1.765 4.165 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 3.470 2.430 4.165 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.545 2.120 3.045 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.470 3.650 4.165 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.410 2.630 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.980 0.520 3.860 ;
        RECT  0.120 0.845 0.520 1.185 ;
        RECT  0.120 0.845 0.410 3.860 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 3.470 5.125 4.000 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.880 3.470 4.165 5.280 ;
        RECT  0.900 3.020 1.220 3.345 ;
        RECT  0.900 3.020 1.185 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  0.940 -0.400 1.860 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.940 1.460 3.920 1.800 ;
        RECT  0.940 1.460 1.280 1.995 ;
        RECT  4.380 1.360 5.490 1.700 ;
        RECT  0.640 2.350 1.855 2.690 ;
        RECT  1.555 2.350 1.855 3.240 ;
        RECT  5.210 1.360 5.490 3.240 ;
        RECT  1.555 2.900 5.490 3.240 ;
        RECT  3.620 0.710 5.490 1.060 ;
        RECT  0.940 1.460 2.40 1.800 ;
        RECT  1.555 2.900 4.40 3.240 ;
    END
END OA222X1

MACRO OA222X0
    CLASS CORE ;
    FOREIGN OA222X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.060 2.250 1.765 2.630 ;
        RECT  1.060 2.135 1.400 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.730 3.470 2.395 3.865 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.300 2.250 3.025 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 3.465 3.660 3.820 ;
        RECT  2.965 3.465 3.270 3.825 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.510 ;
        RECT  0.125 2.815 0.520 3.130 ;
        RECT  0.125 1.030 0.520 1.510 ;
        RECT  0.125 1.030 0.355 3.130 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.240 3.470 4.915 3.865 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.570 2.230 4.285 2.630 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.290 4.055 3.630 5.280 ;
        RECT  3.320 4.050 3.630 5.280 ;
        RECT  0.780 3.985 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  1.245 -0.400 1.585 1.845 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.735 0.715 3.785 1.055 ;
        RECT  2.735 0.715 3.075 1.845 ;
        RECT  4.135 1.210 4.860 1.550 ;
        RECT  4.520 2.815 4.860 3.155 ;
        RECT  4.630 1.210 4.860 3.155 ;
        RECT  0.925 2.870 4.860 3.155 ;
        RECT  0.925 2.870 1.155 3.755 ;
        RECT  0.460 3.450 1.155 3.755 ;
        RECT  0.925 2.870 3.30 3.155 ;
    END
END OA222X0

MACRO OA221X4
    CLASS CORE ;
    FOREIGN OA221X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.580 2.100 3.045 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.880 2.055 4.305 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.055 5.565 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.120 6.280 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.055 4.935 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.450 3.320 1.960 4.160 ;
        RECT  1.440 1.290 1.840 1.630 ;
        RECT  1.450 1.290 1.680 4.160 ;
        RECT  0.180 2.250 1.680 2.630 ;
        RECT  1.440 1.290 1.680 2.630 ;
        RECT  0.180 0.700 0.520 4.160 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 3.320 6.030 5.280 ;
        RECT  2.340 3.320 3.355 5.280 ;
        RECT  0.900 2.910 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  3.580 -0.400 3.920 0.710 ;
        RECT  2.060 -0.400 2.400 0.710 ;
        RECT  0.940 -0.400 1.280 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.820 0.820 3.160 1.825 ;
        RECT  4.880 1.280 5.220 1.825 ;
        RECT  2.820 1.595 5.220 1.825 ;
        RECT  4.160 0.820 5.945 1.050 ;
        RECT  4.160 0.820 4.500 1.365 ;
        RECT  5.600 0.820 5.945 1.700 ;
        RECT  6.320 0.820 6.760 1.700 ;
        RECT  1.910 2.390 2.250 3.090 ;
        RECT  1.910 2.860 6.760 3.090 ;
        RECT  4.355 2.860 4.695 4.160 ;
        RECT  6.530 0.820 6.760 4.160 ;
        RECT  6.410 2.860 6.760 4.160 ;
        RECT  2.820 1.595 4.20 1.825 ;
        RECT  1.910 2.860 5.80 3.090 ;
    END
END OA221X4

MACRO OA221X2
    CLASS CORE ;
    FOREIGN OA221X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.940 2.250 2.395 2.750 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.250 3.045 2.750 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.695 2.750 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.925 2.250 4.510 2.685 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 3.105 1.240 4.025 ;
        RECT  0.750 0.820 1.240 1.160 ;
        RECT  0.750 0.820 0.980 4.025 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.470 1.480 4.920 2.020 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.390 3.440 4.730 5.280 ;
        RECT  1.680 3.440 2.020 5.280 ;
        RECT  0.180 3.105 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  1.620 -0.400 2.430 1.160 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.650 1.090 3.990 2.020 ;
        RECT  1.530 1.680 3.990 2.020 ;
        RECT  1.530 1.680 1.870 2.030 ;
        RECT  2.890 0.630 4.775 0.860 ;
        RECT  2.890 0.630 3.230 1.170 ;
        RECT  4.425 0.630 4.775 1.170 ;
        RECT  1.270 2.350 1.700 2.690 ;
        RECT  1.470 2.350 1.700 3.210 ;
        RECT  1.470 2.980 5.500 3.210 ;
        RECT  3.045 2.980 3.385 4.025 ;
        RECT  5.150 0.830 5.500 4.025 ;
        RECT  1.530 1.680 2.80 2.020 ;
        RECT  1.470 2.980 4.80 3.210 ;
    END
END OA221X2

MACRO OA221X1
    CLASS CORE ;
    FOREIGN OA221X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 3.470 1.765 4.165 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 3.470 2.430 4.165 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.545 2.120 3.045 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.060 3.675 2.670 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.030 4.320 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.980 0.520 3.850 ;
        RECT  0.120 0.850 0.520 1.190 ;
        RECT  0.120 0.850 0.410 3.850 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  0.940 -0.400 1.860 0.940 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.760 3.470 4.100 5.280 ;
        RECT  0.900 3.020 1.220 3.345 ;
        RECT  0.900 3.020 1.185 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.940 1.460 3.920 1.800 ;
        RECT  0.940 1.460 1.280 1.995 ;
        RECT  4.340 0.700 4.860 1.040 ;
        RECT  0.640 2.350 1.855 2.690 ;
        RECT  1.555 2.350 1.855 3.240 ;
        RECT  4.575 0.700 4.860 3.240 ;
        RECT  1.555 2.900 4.860 3.240 ;
        RECT  0.940 1.460 2.30 1.800 ;
        RECT  1.555 2.900 3.70 3.240 ;
    END
END OA221X1

MACRO OA221X0
    CLASS CORE ;
    FOREIGN OA221X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.225 1.400 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.520 2.070 3.875 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.235 2.585 2.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.815 0.630 3.485 1.020 ;
        RECT  2.815 2.425 3.255 2.765 ;
        RECT  2.815 0.630 3.045 2.765 ;
        RECT  2.645 1.030 3.045 1.410 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.170 0.785 1.510 ;
        RECT  0.125 3.005 0.520 3.320 ;
        RECT  0.125 1.030 0.520 1.510 ;
        RECT  0.125 1.030 0.355 3.320 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.945 1.030 4.285 2.005 ;
        RECT  3.905 1.030 4.285 1.410 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.050 4.170 3.390 5.280 ;
        RECT  0.780 4.185 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.245 -0.400 1.585 1.845 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.385 1.250 3.675 1.765 ;
        RECT  0.925 3.005 2.530 3.290 ;
        RECT  3.485 1.555 3.715 3.775 ;
        RECT  2.300 3.005 2.530 3.775 ;
        RECT  3.485 3.435 4.190 3.775 ;
        RECT  2.300 3.490 4.190 3.775 ;
        RECT  0.925 3.005 1.155 3.955 ;
        RECT  0.460 3.640 1.155 3.955 ;
    END
END OA221X0

MACRO OA21X4
    CLASS CORE ;
    FOREIGN OA21X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.140 3.215 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.615 3.840 1.960 4.180 ;
        RECT  1.615 1.280 1.960 1.620 ;
        RECT  1.615 2.955 1.955 4.180 ;
        RECT  1.615 1.280 1.845 4.180 ;
        RECT  0.125 2.400 1.845 2.630 ;
        RECT  0.125 0.700 0.520 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.895 2.140 5.545 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.140 4.515 2.630 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.655 -0.400 3.995 0.990 ;
        RECT  2.195 -0.400 2.535 0.710 ;
        RECT  0.900 -0.400 1.240 1.620 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.135 2.860 5.475 5.280 ;
        RECT  2.340 3.320 3.480 5.280 ;
        RECT  0.900 2.930 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.895 0.820 3.235 1.450 ;
        RECT  4.415 0.820 4.755 1.450 ;
        RECT  2.895 1.220 4.755 1.450 ;
        RECT  5.135 0.820 5.475 1.910 ;
        RECT  3.445 1.680 5.475 1.910 ;
        RECT  2.075 2.410 2.415 2.750 ;
        RECT  2.185 2.410 2.415 3.090 ;
        RECT  3.445 1.680 3.675 3.090 ;
        RECT  2.185 2.860 4.755 3.090 ;
        RECT  4.415 2.860 4.755 4.180 ;
        RECT  3.445 1.680 4.30 1.910 ;
        RECT  2.185 2.860 3.70 3.090 ;
    END
END OA21X4

MACRO OA21X2
    CLASS CORE ;
    FOREIGN OA21X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.955 2.230 2.565 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.750 1.245 3.850 ;
        RECT  0.750 1.240 1.090 3.850 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.650 2.230 4.285 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.470 3.100 4.190 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  2.570 -0.400 2.910 1.540 ;
        RECT  1.310 -0.400 1.650 0.720 ;
        RECT  0.190 -0.400 0.530 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.890 2.860 4.230 5.280 ;
        RECT  1.735 2.860 2.080 5.280 ;
        RECT  0.180 2.750 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.890 1.270 4.230 2.000 ;
        RECT  1.385 1.770 4.230 2.000 ;
        RECT  1.385 1.770 1.725 2.220 ;
        RECT  3.080 1.770 3.420 3.240 ;
        RECT  1.385 1.770 3.10 2.000 ;
    END
END OA21X2

MACRO OA21X1
    CLASS CORE ;
    FOREIGN OA21X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 3.470 1.765 4.165 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 3.470 2.395 4.165 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.545 2.120 3.200 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.900 0.520 3.970 ;
        RECT  0.120 1.265 0.520 1.700 ;
        RECT  0.120 1.265 0.350 3.970 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.095 3.470 3.435 5.280 ;
        RECT  0.900 2.720 1.240 3.060 ;
        RECT  0.900 2.720 1.185 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.000 -0.400 2.340 1.700 ;
        RECT  0.740 -0.400 1.095 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.260 0.630 3.665 0.960 ;
        RECT  0.640 1.940 2.030 2.280 ;
        RECT  1.730 1.940 2.030 3.200 ;
        RECT  3.430 0.630 3.665 3.200 ;
        RECT  1.730 2.860 3.665 3.200 ;
    END
END OA21X1

MACRO OA21X0
    CLASS CORE ;
    FOREIGN OA21X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.725 2.250 1.135 2.580 ;
        RECT  0.725 1.770 1.015 2.580 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.680 3.620 2.020 4.050 ;
        RECT  1.385 3.485 1.750 3.850 ;
        RECT  1.385 3.470 1.740 3.850 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.530 2.155 3.035 2.640 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.170 0.785 1.460 ;
        RECT  0.115 3.890 0.520 4.210 ;
        RECT  0.115 1.030 0.520 1.460 ;
        RECT  0.115 1.030 0.345 4.210 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.560 4.170 2.910 5.280 ;
        RECT  0.930 4.170 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.245 -0.400 1.585 1.835 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.070 0.630 2.970 0.970 ;
        RECT  2.070 0.630 2.300 3.390 ;
        RECT  0.580 2.810 2.310 3.100 ;
        RECT  1.970 2.810 2.310 3.390 ;
    END
END OA21X0

MACRO OA211X4
    CLASS CORE ;
    FOREIGN OA211X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.870 2.120 5.545 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.035 6.185 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.254  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 1.130 1.960 4.160 ;
        RECT  0.180 2.250 1.960 2.630 ;
        RECT  0.180 1.130 0.520 4.160 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.195 2.120 3.675 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.461  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.440 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.060 3.320 5.400 5.280 ;
        RECT  3.190 3.320 3.530 5.280 ;
        RECT  2.340 3.320 2.680 5.280 ;
        RECT  0.900 2.910 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 1.700 ;
        RECT  2.340 -0.400 2.680 1.430 ;
        RECT  0.900 -0.400 1.240 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.190 0.820 4.975 1.050 ;
        RECT  3.190 0.820 3.530 1.430 ;
        RECT  4.630 0.820 4.975 1.700 ;
        RECT  3.910 1.280 4.250 1.890 ;
        RECT  2.190 1.660 4.250 1.890 ;
        RECT  2.190 1.660 2.530 3.090 ;
        RECT  2.190 2.860 6.120 3.090 ;
        RECT  4.340 2.860 4.680 4.160 ;
        RECT  5.780 2.860 6.120 4.160 ;
        RECT  2.190 1.660 3.30 1.890 ;
        RECT  2.190 2.860 5.20 3.090 ;
    END
END OA211X4

MACRO OA211X2
    CLASS CORE ;
    FOREIGN OA211X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.650 1.150 3.560 ;
        RECT  0.755 1.240 1.150 1.580 ;
        RECT  0.755 1.240 1.060 3.560 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.045 3.470 2.395 4.165 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 3.470 3.025 4.165 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.120 3.950 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.360 1.995 4.915 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.760 3.430 4.100 5.280 ;
        RECT  1.530 2.640 1.870 2.980 ;
        RECT  1.530 2.640 1.815 5.280 ;
        RECT  0.250 4.015 0.590 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.520 -0.400 4.860 1.610 ;
        RECT  1.370 -0.400 1.710 0.720 ;
        RECT  0.250 -0.400 0.590 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.700 1.270 3.040 2.280 ;
        RECT  1.290 1.940 3.040 2.280 ;
        RECT  2.810 1.270 3.040 3.200 ;
        RECT  2.810 2.860 4.860 3.200 ;
        RECT  2.810 2.860 3.80 3.200 ;
    END
END OA211X2

MACRO OA211X1
    CLASS CORE ;
    FOREIGN OA211X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.650 0.520 3.970 ;
        RECT  0.120 1.265 0.520 1.700 ;
        RECT  0.120 1.265 0.350 3.970 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 3.470 1.765 4.165 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 3.470 2.395 4.165 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.120 3.320 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.730 1.995 4.285 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.130 3.470 3.470 5.280 ;
        RECT  0.900 2.720 1.240 3.060 ;
        RECT  0.900 2.720 1.185 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.890 -0.400 4.230 1.700 ;
        RECT  0.805 -0.400 1.160 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.070 1.360 2.410 2.280 ;
        RECT  0.640 1.940 2.410 2.280 ;
        RECT  2.110 1.360 2.410 3.200 ;
        RECT  2.110 2.860 4.230 3.200 ;
        RECT  2.110 2.860 3.60 3.200 ;
    END
END OA211X1

MACRO OA211X0
    CLASS CORE ;
    FOREIGN OA211X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.135 1.765 2.630 ;
        RECT  0.725 2.135 1.765 2.365 ;
        RECT  0.725 1.770 1.015 2.365 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.680 3.710 3.025 3.940 ;
        RECT  2.645 3.470 3.025 3.940 ;
        RECT  1.680 3.710 2.020 4.050 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.030 2.765 1.410 ;
        RECT  2.365 0.630 2.765 1.410 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.586  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.170 0.785 1.510 ;
        RECT  0.115 3.470 0.520 4.250 ;
        RECT  0.115 1.170 0.345 4.250 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.040 2.250 3.655 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.560 4.170 2.900 5.280 ;
        RECT  0.930 4.170 1.270 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.260 -0.400 3.600 1.700 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.245 1.495 1.585 1.900 ;
        RECT  1.245 1.670 2.225 1.900 ;
        RECT  0.580 2.595 0.965 2.925 ;
        RECT  0.735 2.595 0.965 3.240 ;
        RECT  1.995 1.670 2.225 3.445 ;
        RECT  0.735 3.010 3.490 3.240 ;
        RECT  1.960 3.010 2.300 3.445 ;
        RECT  3.260 3.010 3.490 4.185 ;
        RECT  3.260 3.845 3.600 4.185 ;
        RECT  0.735 3.010 2.60 3.240 ;
    END
END OA211X0

MACRO NO8X1
    CLASS CORE ;
    FOREIGN NO8X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.385 2.120 8.875 2.460 ;
        RECT  8.315 2.860 8.695 3.240 ;
        RECT  8.385 2.120 8.695 3.240 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.540 4.970 1.770 ;
        RECT  4.630 1.170 4.970 1.770 ;
        RECT  3.905 2.960 4.450 3.880 ;
        RECT  3.905 1.540 4.185 3.880 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.145 3.470 3.675 4.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.720 1.795 3.115 2.135 ;
        RECT  2.720 1.030 3.025 2.135 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.005 1.765 3.240 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.685 2.435 2.320 ;
        END
    END E
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.870 1.670 8.155 2.475 ;
        RECT  7.685 2.245 8.065 2.650 ;
        END
    END G
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.190 1.620 7.530 1.945 ;
        RECT  6.425 1.620 7.530 1.850 ;
        RECT  6.425 1.030 6.805 1.850 ;
        END
    END H
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 1.690 1.135 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.270 3.795 7.610 5.280 ;
        RECT  4.870 2.685 6.050 3.025 ;
        RECT  4.870 2.685 5.210 5.280 ;
        RECT  1.995 3.040 2.325 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  6.990 -0.400 8.530 0.710 ;
        RECT  2.630 -0.400 3.940 0.745 ;
        RECT  0.980 -0.400 1.320 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.170 1.170 2.120 1.455 ;
        RECT  0.170 1.170 0.520 1.510 ;
        RECT  0.170 1.170 0.470 4.250 ;
        RECT  0.170 3.165 0.705 3.505 ;
        RECT  0.170 3.165 0.510 4.250 ;
        RECT  4.170 0.630 5.320 0.915 ;
        RECT  4.170 0.630 4.400 1.310 ;
        RECT  3.255 1.080 4.400 1.310 ;
        RECT  3.255 1.080 3.575 1.530 ;
        RECT  3.345 1.080 3.575 3.240 ;
        RECT  3.210 2.955 3.575 3.240 ;
        RECT  5.330 1.170 5.670 2.335 ;
        RECT  4.415 2.000 5.670 2.335 ;
        RECT  4.415 2.105 6.810 2.335 ;
        RECT  6.470 2.105 6.810 3.845 ;
        RECT  5.630 3.505 6.810 3.845 ;
        RECT  8.930 0.630 9.335 1.395 ;
        RECT  7.590 1.070 9.335 1.395 ;
        RECT  9.105 0.630 9.335 3.200 ;
        RECT  8.930 2.860 9.160 4.250 ;
        RECT  7.840 3.945 9.160 4.250 ;
        RECT  4.415 2.105 5.90 2.335 ;
    END
END NO8X1

MACRO NO8X0
    CLASS CORE ;
    FOREIGN NO8X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.645 7.580 1.930 ;
        RECT  6.425 1.030 6.805 1.930 ;
        END
    END H
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 1.690 1.135 2.380 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.690 2.435 2.325 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.525 2.090 8.875 2.430 ;
        RECT  8.315 2.865 8.755 3.250 ;
        RECT  8.525 2.090 8.755 3.250 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.250 8.260 2.640 ;
        RECT  7.920 1.670 8.260 2.640 ;
        END
    END G
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.745 3.120 2.030 ;
        RECT  2.780 1.695 3.115 2.030 ;
        RECT  2.780 1.030 3.025 2.030 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.090 1.765 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.408  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.330 1.540 4.970 1.820 ;
        RECT  4.630 1.170 4.970 1.820 ;
        RECT  3.955 3.270 4.560 3.610 ;
        RECT  4.330 1.540 4.560 3.610 ;
        RECT  3.955 3.270 4.285 3.850 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.220 3.725 3.850 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  6.990 -0.400 8.530 0.710 ;
        RECT  2.630 -0.400 3.940 0.745 ;
        RECT  0.980 -0.400 1.320 0.995 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.410 3.290 7.750 5.280 ;
        RECT  4.940 2.620 6.080 2.910 ;
        RECT  4.940 2.620 5.280 5.280 ;
        RECT  2.500 2.620 2.845 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.780 1.170 2.120 1.460 ;
        RECT  0.180 1.225 2.120 1.460 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  0.180 1.170 0.410 3.325 ;
        RECT  0.180 3.040 1.145 3.325 ;
        RECT  0.690 3.040 1.145 3.380 ;
        RECT  0.690 3.040 1.030 3.905 ;
        RECT  4.170 0.630 5.120 0.915 ;
        RECT  4.170 0.630 4.400 1.310 ;
        RECT  3.255 1.080 4.400 1.310 ;
        RECT  3.255 1.080 4.070 1.510 ;
        RECT  3.730 1.080 4.070 2.870 ;
        RECT  5.330 1.095 5.670 2.390 ;
        RECT  4.790 2.050 5.670 2.390 ;
        RECT  4.790 2.160 6.880 2.390 ;
        RECT  6.540 2.160 6.880 3.610 ;
        RECT  5.740 3.270 6.880 3.610 ;
        RECT  8.890 0.630 9.335 1.390 ;
        RECT  7.590 1.070 9.335 1.390 ;
        RECT  9.105 0.630 9.335 2.980 ;
        RECT  8.985 2.640 9.215 3.910 ;
        RECT  7.995 3.570 9.215 3.910 ;
        RECT  4.790 2.160 5.80 2.390 ;
    END
END NO8X0

MACRO NO7X1
    CLASS CORE ;
    FOREIGN NO7X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.685 2.435 2.320 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 1.850 1.135 2.630 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.145 3.470 3.665 4.100 ;
        END
    END A
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.280 1.615 7.620 1.930 ;
        RECT  6.425 1.615 7.620 1.845 ;
        RECT  6.425 1.030 6.805 1.845 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.000 1.765 3.240 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.720 1.795 3.115 2.135 ;
        RECT  2.720 1.030 3.025 2.135 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.815  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.245 1.540 4.970 1.770 ;
        RECT  4.630 1.170 4.970 1.770 ;
        RECT  3.905 3.460 4.475 3.880 ;
        RECT  4.245 1.540 4.475 3.880 ;
        RECT  4.095 2.960 4.475 3.880 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.960 1.670 8.245 2.480 ;
        RECT  7.685 2.250 8.065 2.640 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.990 -0.400 8.530 0.710 ;
        RECT  2.630 -0.400 3.940 0.745 ;
        RECT  0.980 -0.400 1.320 0.995 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.270 3.660 7.610 5.280 ;
        RECT  4.870 2.690 6.130 3.030 ;
        RECT  4.870 2.690 5.210 5.280 ;
        RECT  2.035 3.120 2.365 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.780 1.170 2.120 1.455 ;
        RECT  0.170 1.225 2.120 1.455 ;
        RECT  0.170 1.170 0.520 1.510 ;
        RECT  0.170 1.170 0.410 4.250 ;
        RECT  0.170 3.190 0.745 3.530 ;
        RECT  0.170 3.190 0.510 4.250 ;
        RECT  4.170 0.630 5.320 0.915 ;
        RECT  4.170 0.630 4.400 1.310 ;
        RECT  3.255 1.080 4.400 1.310 ;
        RECT  3.255 1.080 3.575 1.530 ;
        RECT  3.345 1.080 3.575 3.240 ;
        RECT  3.210 2.955 3.575 3.240 ;
        RECT  5.330 1.170 5.670 2.335 ;
        RECT  4.705 2.000 5.670 2.335 ;
        RECT  4.705 2.105 6.850 2.335 ;
        RECT  6.510 2.105 6.850 3.830 ;
        RECT  5.630 3.490 6.850 3.830 ;
        RECT  7.590 1.070 8.705 1.385 ;
        RECT  8.475 1.070 8.705 3.115 ;
        RECT  8.260 2.775 8.490 4.250 ;
        RECT  7.840 3.910 8.490 4.250 ;
        RECT  4.705 2.105 5.20 2.335 ;
    END
END NO7X1

MACRO NO7X0
    CLASS CORE ;
    FOREIGN NO7X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 2.030 1.135 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.685 2.435 2.320 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.960 1.670 8.245 2.495 ;
        RECT  7.685 2.250 8.065 2.630 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.280 1.615 7.620 1.930 ;
        RECT  6.425 1.615 7.620 1.875 ;
        RECT  6.425 1.030 6.805 1.875 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.090 1.765 3.240 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.745 3.120 2.030 ;
        RECT  2.780 1.695 3.115 2.030 ;
        RECT  2.780 1.030 3.025 2.030 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.175 3.725 3.850 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.408  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.245 1.540 4.970 1.770 ;
        RECT  4.630 1.170 4.970 1.770 ;
        RECT  3.955 3.230 4.475 3.850 ;
        RECT  4.245 1.540 4.475 3.850 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.990 -0.400 8.530 0.710 ;
        RECT  2.630 -0.400 3.940 0.745 ;
        RECT  0.980 -0.400 1.320 0.995 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.270 3.380 7.610 5.280 ;
        RECT  4.870 2.565 6.010 2.870 ;
        RECT  4.870 2.565 5.210 5.280 ;
        RECT  2.500 2.620 2.845 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  1.780 1.170 2.120 1.455 ;
        RECT  0.180 1.225 2.120 1.455 ;
        RECT  0.180 1.225 1.770 1.510 ;
        RECT  0.180 1.170 0.410 3.325 ;
        RECT  0.180 3.040 1.145 3.325 ;
        RECT  0.690 3.040 1.145 3.380 ;
        RECT  0.690 3.040 1.030 3.905 ;
        RECT  4.170 0.630 5.120 0.915 ;
        RECT  4.170 0.630 4.400 1.310 ;
        RECT  3.255 1.080 4.400 1.310 ;
        RECT  3.255 1.080 4.015 1.510 ;
        RECT  3.730 1.080 4.015 2.870 ;
        RECT  5.330 1.095 5.670 2.335 ;
        RECT  4.705 2.000 5.670 2.335 ;
        RECT  4.705 2.105 6.810 2.335 ;
        RECT  6.470 2.105 6.810 3.570 ;
        RECT  5.670 3.230 6.810 3.570 ;
        RECT  7.590 1.070 8.705 1.385 ;
        RECT  8.475 1.070 8.705 3.070 ;
        RECT  8.300 2.730 8.530 4.000 ;
        RECT  7.840 3.660 8.530 4.000 ;
        RECT  4.705 2.105 5.80 2.335 ;
    END
END NO7X0

MACRO NO6X4
    CLASS CORE ;
    FOREIGN NO6X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.860 1.135 3.240 ;
        RECT  0.750 2.135 0.980 3.240 ;
        RECT  0.575 2.135 0.980 2.480 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.100 3.045 2.625 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 1.040 9.275 4.160 ;
        RECT  7.730 2.205 9.275 2.655 ;
        RECT  7.490 3.115 7.960 4.160 ;
        RECT  7.730 1.040 7.960 4.160 ;
        RECT  7.490 1.040 7.960 1.380 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 2.250 1.765 2.625 ;
        RECT  1.210 1.780 1.520 2.625 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.140 3.675 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.140 4.400 2.630 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 1.720 2.400 2.030 ;
        RECT  1.915 1.640 2.400 2.030 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.210 -0.400 8.550 1.510 ;
        RECT  6.730 -0.400 7.070 1.000 ;
        RECT  3.780 -0.400 4.120 0.710 ;
        RECT  2.380 -0.400 2.720 0.710 ;
        RECT  0.900 -0.400 1.240 1.090 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.210 2.920 8.550 5.280 ;
        RECT  6.770 3.180 7.110 5.280 ;
        RECT  5.330 2.720 5.670 5.280 ;
        RECT  1.960 2.855 2.770 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.150 1.400 4.890 1.715 ;
        RECT  4.640 1.400 4.890 2.490 ;
        RECT  4.640 2.150 6.150 2.490 ;
        RECT  4.640 1.400 4.880 3.090 ;
        RECT  4.290 2.860 4.640 4.175 ;
        RECT  1.470 0.940 5.350 1.170 ;
        RECT  1.470 0.940 1.960 1.280 ;
        RECT  0.115 0.785 0.520 1.550 ;
        RECT  1.470 0.940 1.700 1.550 ;
        RECT  0.115 1.320 1.700 1.550 ;
        RECT  5.120 0.940 5.350 1.920 ;
        RECT  5.120 1.690 6.720 1.920 ;
        RECT  6.490 1.690 6.720 2.490 ;
        RECT  6.490 2.150 6.825 2.490 ;
        RECT  0.115 0.785 0.345 4.175 ;
        RECT  0.115 2.715 0.520 4.175 ;
        RECT  5.580 0.700 5.920 1.460 ;
        RECT  5.580 1.230 7.260 1.460 ;
        RECT  7.030 1.230 7.260 2.040 ;
        RECT  7.055 1.890 7.500 2.230 ;
        RECT  7.055 1.890 7.320 2.950 ;
        RECT  6.050 2.720 7.320 2.950 ;
        RECT  6.050 2.720 6.390 4.180 ;
        RECT  1.470 0.940 4.30 1.170 ;
    END
END NO6X4

MACRO NO6X2
    CLASS CORE ;
    FOREIGN NO6X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.785 2.300 6.355 2.700 ;
        RECT  5.785 2.250 6.200 2.700 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.590 2.120 1.085 2.685 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.670 2.050 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.640 6.985 2.050 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.375 2.250 4.925 2.630 ;
        RECT  4.330 3.040 4.670 3.960 ;
        RECT  4.375 2.250 4.670 3.960 ;
        RECT  4.375 1.680 4.605 3.960 ;
        RECT  4.230 1.680 4.605 2.020 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 2.250 2.440 2.685 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.315 2.320 1.715 3.240 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.105 2.960 5.445 5.280 ;
        RECT  3.610 3.080 3.950 5.280 ;
        RECT  2.170 3.040 2.510 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.410 -0.400 6.750 0.710 ;
        RECT  4.890 -0.400 5.230 0.950 ;
        RECT  2.340 -0.400 2.680 1.430 ;
        RECT  0.900 -0.400 1.240 1.430 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.180 0.520 1.890 ;
        RECT  1.620 1.180 1.960 1.890 ;
        RECT  0.115 1.660 2.900 1.890 ;
        RECT  2.575 1.660 2.900 2.060 ;
        RECT  0.115 1.180 0.360 3.330 ;
        RECT  0.350 2.990 0.690 3.955 ;
        RECT  3.130 0.700 3.870 0.990 ;
        RECT  3.130 0.700 3.360 2.850 ;
        RECT  3.130 2.520 4.145 2.850 ;
        RECT  2.890 2.635 3.230 3.960 ;
        RECT  5.650 1.100 5.990 1.410 ;
        RECT  4.745 1.180 7.445 1.410 ;
        RECT  7.040 1.110 7.445 1.410 ;
        RECT  3.590 1.220 4.935 1.450 ;
        RECT  3.590 1.220 3.930 2.150 ;
        RECT  7.215 1.110 7.445 3.205 ;
        RECT  6.925 2.975 7.265 4.080 ;
        RECT  0.115 1.660 1.70 1.890 ;
        RECT  4.745 1.180 6.30 1.410 ;
    END
END NO6X2

MACRO NO6X1
    CLASS CORE ;
    FOREIGN NO6X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.700 1.690 1.135 2.375 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.620 5.640 1.930 ;
        RECT  4.535 1.030 4.915 1.930 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.980 1.670 6.320 2.010 ;
        RECT  5.795 2.250 6.260 2.650 ;
        RECT  5.980 1.670 6.260 2.650 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.690 2.435 2.320 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 1.690 1.765 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.870 1.030 3.655 1.485 ;
        RECT  3.090 2.335 3.430 3.550 ;
        RECT  2.870 1.030 3.100 2.565 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.635 2.105 6.985 2.445 ;
        RECT  6.425 2.860 6.865 3.250 ;
        RECT  6.635 2.105 6.865 3.250 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.360 2.890 5.700 5.280 ;
        RECT  3.840 2.640 4.180 5.280 ;
        RECT  2.310 2.855 2.650 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.100 -0.400 6.640 0.710 ;
        RECT  0.980 -0.400 2.690 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 1.995 1.460 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  0.180 1.170 0.410 3.110 ;
        RECT  0.180 2.825 1.070 3.110 ;
        RECT  0.540 2.825 1.070 3.165 ;
        RECT  0.540 2.825 0.880 3.960 ;
        RECT  3.885 1.070 4.220 2.030 ;
        RECT  3.330 1.715 4.220 2.030 ;
        RECT  3.935 1.070 4.220 2.390 ;
        RECT  3.935 2.160 4.940 2.390 ;
        RECT  4.600 2.160 4.940 2.980 ;
        RECT  7.000 0.630 7.445 1.395 ;
        RECT  5.700 1.070 7.445 1.395 ;
        RECT  7.215 0.630 7.445 3.215 ;
        RECT  7.095 2.875 7.325 4.250 ;
        RECT  6.105 3.955 7.325 4.250 ;
    END
END NO6X1

MACRO NO6X0
    CLASS CORE ;
    FOREIGN NO6X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.640 0.505 2.265 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 1.635 5.060 2.040 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.250 5.740 2.630 ;
        RECT  5.400 1.690 5.740 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.970 2.080 6.355 2.420 ;
        RECT  5.795 2.860 6.200 3.240 ;
        RECT  5.970 2.080 6.200 3.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 1.640 2.395 2.100 ;
        RECT  1.855 1.640 2.395 2.035 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.200 2.250 1.765 2.630 ;
        RECT  1.200 1.690 1.540 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.562  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 0.630 3.120 1.410 ;
        RECT  2.620 2.640 2.960 2.980 ;
        RECT  2.625 0.630 2.855 2.980 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.890 3.360 5.230 5.280 ;
        RECT  3.220 3.380 3.560 5.280 ;
        RECT  1.840 2.925 2.180 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.510 -0.400 6.050 0.710 ;
        RECT  0.880 -0.400 2.395 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.090 1.820 1.410 ;
        RECT  0.735 1.090 1.805 1.415 ;
        RECT  0.735 1.090 0.965 2.870 ;
        RECT  0.180 2.640 0.965 2.870 ;
        RECT  0.180 2.640 0.520 3.890 ;
        RECT  3.480 0.630 3.820 2.390 ;
        RECT  3.085 2.050 3.820 2.390 ;
        RECT  3.085 2.160 4.250 2.390 ;
        RECT  4.020 2.160 4.250 3.050 ;
        RECT  4.020 2.710 4.360 3.050 ;
        RECT  6.410 0.630 6.815 1.410 ;
        RECT  5.110 1.070 6.815 1.410 ;
        RECT  6.585 0.630 6.815 3.050 ;
        RECT  6.430 2.710 6.660 3.980 ;
        RECT  5.475 3.640 6.660 3.980 ;
    END
END NO6X0

MACRO NO6I5X4
    CLASS CORE ;
    FOREIGN NO6I5X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 3.430 3.130 3.930 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.230 2.120 3.710 2.635 ;
        RECT  3.220 2.120 3.710 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.215  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.000 3.105 9.340 3.895 ;
        RECT  9.000 3.095 9.330 3.895 ;
        RECT  9.000 2.490 9.230 3.895 ;
        RECT  7.430 1.405 9.090 1.690 ;
        RECT  7.560 2.490 9.230 2.720 ;
        RECT  8.315 1.405 8.695 2.720 ;
        RECT  7.560 2.490 7.900 3.895 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.880 2.395 3.240 ;
        RECT  1.995 1.880 2.395 2.220 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 2.210 1.765 2.650 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.460 3.235 11.845 3.850 ;
        RECT  11.260 3.235 11.845 3.575 ;
        END
    END EN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.620 1.030 11.215 1.410 ;
        RECT  10.620 0.630 10.850 1.410 ;
        RECT  10.330 0.630 10.850 0.940 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.890 3.805 11.230 5.280 ;
        RECT  8.280 2.950 8.620 5.280 ;
        RECT  6.840 2.910 7.180 5.280 ;
        RECT  5.400 3.150 5.740 5.280 ;
        RECT  3.380 3.650 3.720 5.280 ;
        RECT  2.060 3.650 2.400 5.280 ;
        RECT  0.740 4.150 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  11.080 -0.400 11.425 0.800 ;
        RECT  9.490 -0.400 9.830 0.715 ;
        RECT  8.190 -0.400 8.530 0.710 ;
        RECT  6.575 -0.400 6.915 0.710 ;
        RECT  3.170 -0.400 3.455 0.785 ;
        RECT  0.940 -0.400 1.280 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.240 0.520 1.580 ;
        RECT  0.130 1.240 0.360 3.750 ;
        RECT  0.130 2.830 0.520 3.750 ;
        RECT  0.130 3.520 1.650 3.750 ;
        RECT  1.310 3.520 1.650 4.250 ;
        RECT  1.770 0.640 2.110 1.440 ;
        RECT  0.750 1.210 2.110 1.440 ;
        RECT  0.590 2.260 0.980 2.600 ;
        RECT  0.750 1.210 0.980 3.220 ;
        RECT  0.750 2.880 1.785 3.220 ;
        RECT  3.685 0.630 4.160 0.940 ;
        RECT  2.470 0.640 2.810 1.245 ;
        RECT  3.685 0.630 3.915 1.245 ;
        RECT  2.470 1.015 3.915 1.245 ;
        RECT  2.760 1.015 2.990 3.195 ;
        RECT  2.760 2.855 3.160 3.195 ;
        RECT  4.115 1.360 4.480 1.700 ;
        RECT  4.090 1.395 4.480 1.700 ;
        RECT  4.250 2.120 5.885 2.350 ;
        RECT  5.600 2.120 5.885 2.460 ;
        RECT  4.250 1.360 4.480 3.170 ;
        RECT  4.140 2.830 4.480 3.170 ;
        RECT  4.760 0.700 5.100 1.700 ;
        RECT  4.760 1.470 6.345 1.700 ;
        RECT  7.100 1.920 7.530 2.260 ;
        RECT  7.100 1.920 7.330 2.680 ;
        RECT  6.115 2.450 7.330 2.680 ;
        RECT  6.115 1.470 6.345 2.920 ;
        RECT  4.790 2.690 6.460 2.920 ;
        RECT  4.790 2.690 5.020 3.845 ;
        RECT  4.680 3.505 5.020 3.845 ;
        RECT  6.120 2.450 6.460 4.160 ;
        RECT  6.575 0.945 9.710 1.175 ;
        RECT  9.480 1.240 10.390 1.580 ;
        RECT  6.575 0.945 6.860 2.220 ;
        RECT  9.480 0.945 9.710 2.920 ;
        RECT  9.700 2.690 10.040 3.960 ;
        RECT  9.940 2.120 11.790 2.460 ;
        RECT  11.450 1.340 11.790 3.005 ;
        RECT  6.575 0.945 8.70 1.175 ;
    END
END NO6I5X4

MACRO NO6I5X2
    CLASS CORE ;
    FOREIGN NO6I5X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 3.450 1.830 3.985 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.855 1.345 2.195 ;
        RECT  0.755 1.855 1.135 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.650 1.405 7.880 3.490 ;
        RECT  7.320 3.260 7.660 4.180 ;
        RECT  7.390 1.405 7.880 1.690 ;
        RECT  7.055 3.470 7.660 3.850 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.035 1.695 2.670 2.040 ;
        RECT  2.035 1.635 2.470 2.040 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.270 3.320 2.630 ;
        RECT  2.970 2.120 3.320 2.630 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.000 3.235 10.585 3.850 ;
        END
    END EN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.360 1.030 9.955 1.410 ;
        RECT  9.070 0.780 9.590 1.120 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.430 3.650 9.770 5.280 ;
        RECT  8.040 3.660 8.380 5.280 ;
        RECT  6.560 4.025 6.900 5.280 ;
        RECT  5.280 3.220 5.620 5.280 ;
        RECT  3.460 3.460 3.800 5.280 ;
        RECT  2.060 3.610 2.400 5.280 ;
        RECT  0.740 3.460 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.820 -0.400 10.165 0.800 ;
        RECT  7.990 -0.400 8.330 0.710 ;
        RECT  6.760 -0.400 7.100 0.710 ;
        RECT  3.640 -0.400 3.980 0.780 ;
        RECT  1.160 -0.400 1.500 0.790 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.470 3.935 ;
        RECT  0.180 2.690 0.510 3.935 ;
        RECT  0.460 0.650 0.930 0.940 ;
        RECT  0.700 0.650 0.930 1.250 ;
        RECT  2.010 0.630 2.350 1.250 ;
        RECT  0.700 1.020 2.350 1.250 ;
        RECT  1.575 1.020 1.805 3.005 ;
        RECT  1.495 2.665 1.840 3.005 ;
        RECT  2.635 1.160 3.780 1.465 ;
        RECT  3.550 1.730 4.370 2.070 ;
        RECT  3.550 1.160 3.780 3.130 ;
        RECT  2.760 2.900 3.780 3.130 ;
        RECT  2.760 2.900 3.100 3.800 ;
        RECT  4.440 1.170 4.830 1.510 ;
        RECT  4.600 1.880 5.380 2.220 ;
        RECT  4.600 1.170 4.830 2.530 ;
        RECT  4.020 2.300 4.830 2.530 ;
        RECT  4.020 2.300 4.360 3.020 ;
        RECT  5.140 0.820 5.480 1.650 ;
        RECT  5.140 1.420 5.840 1.650 ;
        RECT  5.610 1.420 5.840 2.990 ;
        RECT  5.610 2.650 7.420 2.990 ;
        RECT  4.630 2.760 7.420 2.990 ;
        RECT  6.000 2.650 6.340 3.555 ;
        RECT  4.630 2.760 4.860 3.750 ;
        RECT  4.520 3.410 4.860 3.750 ;
        RECT  6.480 0.945 8.425 1.175 ;
        RECT  8.195 1.350 9.130 1.690 ;
        RECT  6.480 0.945 6.820 2.235 ;
        RECT  8.195 0.945 8.425 2.970 ;
        RECT  8.195 2.630 8.780 2.970 ;
        RECT  8.655 2.060 10.530 2.400 ;
        RECT  10.190 1.340 10.530 2.980 ;
        RECT  4.630 2.760 6.90 2.990 ;
    END
END NO6I5X2

MACRO NO6I5X1
    CLASS CORE ;
    FOREIGN NO6I5X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 3.450 1.830 3.985 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.855 1.345 2.195 ;
        RECT  0.755 1.855 1.135 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.672  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 3.470 7.440 3.930 ;
        RECT  7.100 1.605 7.330 3.930 ;
        RECT  6.965 1.605 7.330 1.890 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.035 1.700 2.665 2.040 ;
        RECT  2.035 1.640 2.395 2.040 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.270 3.320 2.630 ;
        RECT  2.970 2.130 3.320 2.630 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.470 2.720 9.965 3.190 ;
        END
    END EN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.820 1.030 9.325 1.410 ;
        RECT  8.595 1.690 9.055 2.030 ;
        RECT  8.820 1.030 9.055 2.030 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.720 3.885 9.060 5.280 ;
        RECT  6.305 3.035 6.685 5.280 ;
        RECT  4.860 3.615 5.200 5.280 ;
        RECT  3.460 3.910 3.800 5.280 ;
        RECT  2.060 3.765 2.400 5.280 ;
        RECT  0.740 3.460 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.955 -0.400 9.300 0.785 ;
        RECT  7.360 -0.400 7.700 0.915 ;
        RECT  6.435 -0.400 6.775 0.825 ;
        RECT  3.680 -0.400 4.020 0.710 ;
        RECT  1.155 -0.400 1.495 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.465 3.935 ;
        RECT  0.180 1.220 0.470 3.935 ;
        RECT  0.180 2.690 0.510 3.935 ;
        RECT  0.460 0.650 0.925 0.940 ;
        RECT  2.010 0.630 2.350 0.950 ;
        RECT  0.695 0.940 2.240 1.170 ;
        RECT  1.575 0.940 1.805 3.005 ;
        RECT  1.495 2.665 1.840 3.005 ;
        RECT  2.690 1.160 3.780 1.465 ;
        RECT  3.550 1.750 4.370 2.090 ;
        RECT  3.550 1.160 3.780 3.140 ;
        RECT  2.760 2.910 3.780 3.140 ;
        RECT  2.760 2.910 3.100 3.900 ;
        RECT  4.020 2.640 4.920 2.925 ;
        RECT  4.480 0.720 5.345 1.090 ;
        RECT  4.805 1.470 5.145 2.370 ;
        RECT  4.805 2.140 6.870 2.370 ;
        RECT  5.635 2.140 6.870 2.480 ;
        RECT  4.100 3.155 5.920 3.385 ;
        RECT  4.100 3.155 4.440 3.760 ;
        RECT  5.635 2.140 5.920 3.875 ;
        RECT  5.580 3.155 5.920 3.875 ;
        RECT  5.865 0.630 6.205 1.375 ;
        RECT  8.160 0.720 8.500 1.375 ;
        RECT  5.865 1.145 8.500 1.375 ;
        RECT  7.565 1.145 7.795 3.275 ;
        RECT  7.565 2.935 8.070 3.275 ;
        RECT  9.560 1.160 9.900 2.490 ;
        RECT  8.025 2.260 9.900 2.490 ;
        RECT  8.025 2.260 9.240 2.600 ;
        RECT  9.010 2.260 9.240 3.655 ;
        RECT  9.010 3.420 9.900 3.655 ;
        RECT  9.560 3.420 9.900 3.710 ;
        RECT  4.805 2.140 5.70 2.370 ;
        RECT  5.865 1.145 7.80 1.375 ;
    END
END NO6I5X1

MACRO NO6I5X0
    CLASS CORE ;
    FOREIGN NO6I5X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 3.330 1.845 3.860 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.960 1.345 2.300 ;
        RECT  0.755 1.960 1.135 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.444  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.885 7.420 3.240 ;
        RECT  6.425 2.860 7.250 3.240 ;
        RECT  7.020 1.635 7.250 3.240 ;
        RECT  6.900 1.635 7.250 1.865 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.840 2.220 3.470 2.560 ;
        RECT  2.840 1.030 3.070 2.560 ;
        RECT  2.645 1.030 3.070 1.410 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.035 1.640 2.610 2.065 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.880 3.245 9.325 3.850 ;
        END
    END EN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.940 1.855 8.695 2.195 ;
        RECT  8.315 1.640 8.695 2.195 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.310 3.560 8.650 5.280 ;
        RECT  6.280 3.580 6.620 5.280 ;
        RECT  5.080 3.635 5.420 5.280 ;
        RECT  3.580 3.425 3.920 5.280 ;
        RECT  2.180 3.480 2.520 5.280 ;
        RECT  0.780 3.380 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.130 -0.400 8.470 0.970 ;
        RECT  6.310 -0.400 6.650 0.915 ;
        RECT  4.140 -0.400 4.480 0.710 ;
        RECT  2.510 -0.400 2.850 0.710 ;
        RECT  1.155 -0.400 1.440 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.465 3.830 ;
        RECT  0.180 1.220 0.470 3.830 ;
        RECT  0.180 2.640 0.520 3.830 ;
        RECT  0.460 0.650 0.925 0.940 ;
        RECT  1.810 0.630 2.150 1.170 ;
        RECT  0.695 0.940 2.150 1.170 ;
        RECT  1.575 0.940 1.805 2.930 ;
        RECT  1.575 2.590 1.920 2.930 ;
        RECT  3.340 0.630 3.685 0.960 ;
        RECT  3.455 0.630 3.685 1.940 ;
        RECT  3.455 1.710 4.005 1.940 ;
        RECT  3.700 1.710 4.005 2.050 ;
        RECT  3.700 1.710 3.930 3.095 ;
        RECT  2.880 2.865 3.930 3.095 ;
        RECT  2.880 2.865 3.220 3.690 ;
        RECT  4.140 1.170 4.480 1.510 ;
        RECT  4.235 1.170 4.480 2.940 ;
        RECT  4.235 2.160 5.050 2.445 ;
        RECT  4.235 2.160 4.520 2.940 ;
        RECT  4.180 2.615 4.520 2.940 ;
        RECT  4.840 0.770 5.180 1.930 ;
        RECT  4.840 1.700 5.965 1.930 ;
        RECT  5.680 1.700 5.965 3.405 ;
        RECT  5.680 2.030 6.735 2.370 ;
        RECT  5.680 2.030 6.020 3.405 ;
        RECT  4.280 3.175 6.020 3.405 ;
        RECT  4.280 3.175 4.620 3.750 ;
        RECT  5.740 0.630 6.080 0.915 ;
        RECT  5.850 0.630 6.080 1.375 ;
        RECT  7.330 0.630 7.710 1.375 ;
        RECT  5.850 1.145 7.710 1.375 ;
        RECT  7.480 0.630 7.710 2.655 ;
        RECT  7.650 2.425 7.880 3.930 ;
        RECT  7.080 3.590 7.880 3.930 ;
        RECT  8.910 0.630 9.285 1.510 ;
        RECT  8.965 0.630 9.285 3.015 ;
        RECT  8.910 2.700 9.285 3.015 ;
    END
END NO6I5X0

MACRO NO6I4X4
    CLASS CORE ;
    FOREIGN NO6I4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 3.430 3.130 3.930 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.230 2.120 3.710 2.635 ;
        RECT  3.220 2.120 3.710 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.880 2.640 9.220 3.760 ;
        RECT  7.430 1.405 9.090 1.690 ;
        RECT  7.560 2.640 9.220 2.870 ;
        RECT  8.315 1.405 8.695 2.870 ;
        RECT  7.560 2.640 7.900 3.960 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.880 2.395 3.240 ;
        RECT  1.995 1.880 2.395 2.220 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 2.210 1.765 2.650 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.815 2.120 11.215 3.240 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.240 2.070 10.585 2.640 ;
        RECT  9.910 2.070 10.585 2.410 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 3.470 11.160 5.280 ;
        RECT  8.320 4.160 8.660 5.280 ;
        RECT  6.840 2.910 7.180 5.280 ;
        RECT  5.400 3.150 5.740 5.280 ;
        RECT  3.380 3.650 3.720 5.280 ;
        RECT  2.060 3.650 2.400 5.280 ;
        RECT  0.740 4.150 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.820 -0.400 11.160 1.580 ;
        RECT  9.540 -0.400 9.880 0.715 ;
        RECT  8.190 -0.400 8.530 0.710 ;
        RECT  6.575 -0.400 6.915 0.710 ;
        RECT  3.170 -0.400 3.455 0.785 ;
        RECT  0.940 -0.400 1.280 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.240 0.520 1.580 ;
        RECT  0.130 1.240 0.360 3.750 ;
        RECT  0.130 2.830 0.520 3.750 ;
        RECT  0.130 3.520 1.650 3.750 ;
        RECT  1.310 3.520 1.650 4.250 ;
        RECT  1.770 0.640 2.110 1.440 ;
        RECT  0.750 1.210 2.110 1.440 ;
        RECT  0.590 2.260 0.980 2.600 ;
        RECT  0.750 1.210 0.980 3.220 ;
        RECT  0.750 2.880 1.785 3.220 ;
        RECT  3.685 0.630 4.160 0.940 ;
        RECT  2.470 0.640 2.810 1.245 ;
        RECT  3.685 0.630 3.915 1.245 ;
        RECT  2.470 1.015 3.915 1.245 ;
        RECT  2.760 1.015 2.990 3.195 ;
        RECT  2.760 2.855 3.160 3.195 ;
        RECT  4.115 1.360 4.480 1.700 ;
        RECT  4.090 1.395 4.480 1.700 ;
        RECT  4.140 2.120 5.885 2.350 ;
        RECT  5.600 2.120 5.885 2.460 ;
        RECT  4.140 1.360 4.480 3.170 ;
        RECT  4.760 0.700 5.100 1.700 ;
        RECT  4.760 1.470 6.345 1.700 ;
        RECT  7.100 2.070 7.530 2.410 ;
        RECT  7.100 2.070 7.330 2.680 ;
        RECT  6.115 2.450 7.330 2.680 ;
        RECT  6.115 1.470 6.345 2.920 ;
        RECT  4.790 2.690 6.460 2.920 ;
        RECT  4.790 2.690 5.020 3.845 ;
        RECT  4.680 3.505 5.020 3.845 ;
        RECT  6.120 2.450 6.460 4.160 ;
        RECT  6.575 0.945 9.680 1.175 ;
        RECT  9.450 1.240 10.440 1.580 ;
        RECT  6.575 0.945 6.860 2.220 ;
        RECT  9.450 0.945 9.680 2.920 ;
        RECT  9.670 2.640 10.010 3.960 ;
        RECT  6.575 0.945 8.30 1.175 ;
    END
END NO6I4X4

MACRO NO6I4X2
    CLASS CORE ;
    FOREIGN NO6I4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 3.450 1.830 3.985 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.855 1.345 2.195 ;
        RECT  0.755 1.855 1.135 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.032  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.720 1.405 7.950 3.105 ;
        RECT  7.055 3.470 7.775 3.850 ;
        RECT  7.435 2.870 7.775 3.850 ;
        RECT  7.390 1.405 7.950 1.690 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.035 1.695 2.670 2.040 ;
        RECT  2.035 1.635 2.470 2.040 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.270 3.320 2.630 ;
        RECT  2.970 2.120 3.320 2.630 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 2.060 8.865 2.630 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.555 1.625 9.965 2.225 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.235 2.860 8.575 5.280 ;
        RECT  6.560 4.025 6.900 5.280 ;
        RECT  5.280 3.220 5.620 5.280 ;
        RECT  3.460 3.460 3.800 5.280 ;
        RECT  2.060 3.610 2.400 5.280 ;
        RECT  0.740 3.460 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  9.385 -0.400 9.730 1.040 ;
        RECT  7.990 -0.400 8.330 0.710 ;
        RECT  6.760 -0.400 7.100 0.710 ;
        RECT  3.640 -0.400 3.980 0.780 ;
        RECT  1.160 -0.400 1.500 0.790 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.470 3.935 ;
        RECT  0.180 2.690 0.510 3.935 ;
        RECT  0.460 0.650 0.930 0.940 ;
        RECT  2.010 0.630 2.350 0.950 ;
        RECT  0.700 0.650 0.930 1.250 ;
        RECT  2.010 0.630 2.240 1.250 ;
        RECT  0.700 1.020 2.240 1.250 ;
        RECT  1.575 1.020 1.805 3.005 ;
        RECT  1.495 2.665 1.840 3.005 ;
        RECT  2.635 1.160 3.780 1.465 ;
        RECT  3.550 1.730 4.370 2.070 ;
        RECT  3.550 1.160 3.780 3.230 ;
        RECT  2.760 3.000 3.780 3.230 ;
        RECT  2.760 3.000 3.100 3.800 ;
        RECT  4.440 1.170 4.830 1.510 ;
        RECT  4.600 1.880 5.380 2.220 ;
        RECT  4.600 1.170 4.830 2.530 ;
        RECT  4.020 2.300 4.830 2.530 ;
        RECT  4.020 2.300 4.360 3.020 ;
        RECT  5.140 0.820 5.480 1.650 ;
        RECT  5.140 1.420 6.230 1.650 ;
        RECT  7.050 2.120 7.490 2.460 ;
        RECT  6.000 1.420 6.230 3.555 ;
        RECT  7.050 2.120 7.280 2.695 ;
        RECT  6.000 2.465 7.280 2.695 ;
        RECT  4.630 2.760 6.340 2.990 ;
        RECT  6.000 2.465 6.340 3.555 ;
        RECT  4.630 2.760 4.860 3.750 ;
        RECT  4.520 3.410 4.860 3.750 ;
        RECT  6.590 0.945 9.020 1.175 ;
        RECT  8.790 0.945 9.020 1.690 ;
        RECT  8.790 1.350 9.325 1.690 ;
        RECT  6.590 0.945 6.820 2.235 ;
        RECT  6.480 1.895 6.820 2.235 ;
        RECT  9.095 1.350 9.325 3.200 ;
        RECT  9.095 2.860 9.890 3.200 ;
        RECT  6.590 0.945 8.20 1.175 ;
    END
END NO6I4X2

MACRO NO6I4X1
    CLASS CORE ;
    FOREIGN NO6I4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.495 3.515 8.065 4.010 ;
        END
    END E
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 3.450 1.830 3.985 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.855 1.345 2.195 ;
        RECT  0.755 1.855 1.135 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.670  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.740 2.585 7.350 2.815 ;
        RECT  7.120 1.605 7.350 2.815 ;
        RECT  6.960 1.605 7.350 1.855 ;
        RECT  6.740 3.815 7.080 4.155 ;
        RECT  6.740 2.585 6.970 4.155 ;
        RECT  6.425 2.860 6.970 3.240 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.035 1.680 2.675 2.030 ;
        RECT  2.035 1.630 2.395 2.030 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.260 3.320 2.630 ;
        RECT  2.970 2.120 3.320 2.630 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.165 1.525 8.695 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.295 3.855 8.635 5.280 ;
        RECT  6.005 3.830 6.345 5.280 ;
        RECT  4.860 3.910 5.200 5.280 ;
        RECT  3.460 3.910 3.800 5.280 ;
        RECT  2.060 3.765 2.400 5.280 ;
        RECT  0.740 3.460 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.295 -0.400 8.640 0.735 ;
        RECT  6.410 -0.400 6.750 0.880 ;
        RECT  3.680 -0.400 4.020 0.710 ;
        RECT  1.155 -0.400 1.495 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.465 3.935 ;
        RECT  0.180 1.220 0.470 3.935 ;
        RECT  0.180 2.690 0.510 3.935 ;
        RECT  0.460 0.650 0.925 0.940 ;
        RECT  2.010 0.630 2.350 1.170 ;
        RECT  0.695 0.940 2.350 1.170 ;
        RECT  1.575 0.940 1.805 2.980 ;
        RECT  1.495 2.640 1.840 2.980 ;
        RECT  2.690 1.165 3.780 1.450 ;
        RECT  3.550 1.275 4.540 1.615 ;
        RECT  3.550 1.165 3.780 3.140 ;
        RECT  2.760 2.910 3.780 3.140 ;
        RECT  2.760 2.910 3.100 3.900 ;
        RECT  4.610 2.105 4.950 2.445 ;
        RECT  4.610 2.105 4.840 3.025 ;
        RECT  4.020 2.700 4.840 3.025 ;
        RECT  4.480 0.630 5.340 1.045 ;
        RECT  4.780 1.465 5.120 1.805 ;
        RECT  4.780 1.575 5.705 1.805 ;
        RECT  5.420 1.575 5.705 3.485 ;
        RECT  5.420 2.085 6.890 2.355 ;
        RECT  5.420 2.085 5.760 3.485 ;
        RECT  4.100 3.255 5.760 3.485 ;
        RECT  4.100 3.255 4.440 3.760 ;
        RECT  5.840 0.630 6.180 0.915 ;
        RECT  7.600 0.700 7.940 1.040 ;
        RECT  5.950 0.630 6.180 1.375 ;
        RECT  5.950 1.145 7.840 1.375 ;
        RECT  7.595 1.145 7.840 3.285 ;
        RECT  7.600 0.700 7.840 3.285 ;
        RECT  7.295 3.045 7.840 3.285 ;
    END
END NO6I4X1

MACRO NO6I4X0
    CLASS CORE ;
    FOREIGN NO6I4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 3.335 1.840 3.880 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.345 2.630 ;
        RECT  1.060 1.960 1.345 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.860 7.420 3.240 ;
        RECT  7.020 2.710 7.420 3.240 ;
        RECT  7.020 1.405 7.250 3.240 ;
        RECT  6.900 1.405 7.250 1.745 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.840 2.270 3.470 2.610 ;
        RECT  2.840 1.030 3.070 2.610 ;
        RECT  2.645 1.030 3.070 1.410 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.035 1.640 2.610 2.065 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.650 2.445 8.065 3.240 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.230 1.000 8.695 1.510 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.300 -0.400 8.640 0.710 ;
        RECT  6.230 -0.400 7.040 0.715 ;
        RECT  4.140 -0.400 4.480 0.710 ;
        RECT  2.510 -0.400 2.850 0.710 ;
        RECT  1.155 -0.400 1.450 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.480 3.530 7.410 5.280 ;
        RECT  5.080 3.665 5.420 5.280 ;
        RECT  3.580 3.425 3.920 5.280 ;
        RECT  2.180 3.480 2.520 5.280 ;
        RECT  0.780 3.450 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.465 3.900 ;
        RECT  0.180 1.220 0.470 3.900 ;
        RECT  0.180 2.710 0.520 3.900 ;
        RECT  0.460 0.650 0.925 0.940 ;
        RECT  1.810 0.630 2.150 1.170 ;
        RECT  0.695 0.940 2.150 1.170 ;
        RECT  1.575 0.940 1.805 3.070 ;
        RECT  1.575 2.730 1.920 3.070 ;
        RECT  3.340 0.630 3.685 0.960 ;
        RECT  3.455 0.630 3.685 1.980 ;
        RECT  3.455 1.750 3.985 1.980 ;
        RECT  3.700 1.750 3.985 2.090 ;
        RECT  3.700 1.750 3.930 3.070 ;
        RECT  2.880 2.840 3.930 3.070 ;
        RECT  2.880 2.840 3.220 3.740 ;
        RECT  4.140 1.170 4.480 1.510 ;
        RECT  4.230 1.170 4.480 2.975 ;
        RECT  4.230 2.160 5.050 2.445 ;
        RECT  4.230 2.160 4.520 2.975 ;
        RECT  4.180 2.660 4.520 2.975 ;
        RECT  4.840 0.770 5.180 1.930 ;
        RECT  4.840 1.700 5.965 1.930 ;
        RECT  5.680 1.700 5.965 3.435 ;
        RECT  5.680 1.990 6.790 2.330 ;
        RECT  5.680 1.990 6.020 3.435 ;
        RECT  4.280 3.205 6.020 3.435 ;
        RECT  4.280 3.205 4.620 3.750 ;
        RECT  5.660 0.630 6.000 1.175 ;
        RECT  7.500 0.630 7.840 1.175 ;
        RECT  5.660 0.945 7.840 1.175 ;
        RECT  7.610 0.630 7.840 2.000 ;
        RECT  7.610 1.770 8.640 2.000 ;
        RECT  8.300 1.770 8.640 3.780 ;
        RECT  5.660 0.945 6.80 1.175 ;
    END
END NO6I4X0

MACRO NO6I3X4
    CLASS CORE ;
    FOREIGN NO6I3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.860 1.135 3.240 ;
        RECT  0.575 2.310 0.860 3.240 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.082  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.130 3.585 9.470 4.180 ;
        RECT  8.315 1.345 9.285 1.685 ;
        RECT  7.810 3.585 9.470 3.815 ;
        RECT  7.835 2.660 8.695 2.890 ;
        RECT  8.315 1.345 8.695 2.890 ;
        RECT  7.680 1.345 9.285 1.650 ;
        RECT  7.810 3.430 8.150 3.815 ;
        RECT  7.835 2.660 8.150 3.815 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.230 2.250 1.830 2.650 ;
        RECT  1.190 2.250 1.830 2.635 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.500 1.030 2.395 1.410 ;
        RECT  1.500 0.630 1.840 1.410 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.815 2.120 11.215 3.240 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.240 1.880 10.585 2.640 ;
        RECT  9.975 1.880 10.585 2.220 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.320 2.250 3.780 2.775 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 3.470 11.160 5.280 ;
        RECT  8.370 4.170 8.710 5.280 ;
        RECT  7.250 4.170 7.590 5.280 ;
        RECT  5.730 3.830 6.070 5.280 ;
        RECT  3.280 3.930 3.620 5.280 ;
        RECT  1.990 3.930 2.330 5.280 ;
        RECT  0.880 3.930 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.820 -0.400 11.160 0.715 ;
        RECT  9.700 -0.400 10.040 0.655 ;
        RECT  8.440 -0.400 8.780 0.655 ;
        RECT  6.920 -0.400 7.260 0.655 ;
        RECT  4.420 -0.400 4.760 0.720 ;
        RECT  3.280 -0.400 3.620 0.720 ;
        RECT  2.070 -0.400 2.360 0.800 ;
        RECT  0.980 -0.400 1.270 1.040 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.830 1.500 1.170 2.020 ;
        RECT  0.830 1.790 2.290 2.020 ;
        RECT  2.060 2.260 2.625 2.600 ;
        RECT  2.060 1.790 2.290 3.220 ;
        RECT  1.430 2.880 2.290 3.220 ;
        RECT  0.115 0.700 0.520 1.040 ;
        RECT  4.010 2.310 4.570 2.650 ;
        RECT  0.115 0.700 0.345 4.250 ;
        RECT  4.010 2.310 4.240 3.700 ;
        RECT  0.115 3.470 4.240 3.700 ;
        RECT  0.115 3.470 0.525 4.250 ;
        RECT  2.625 1.375 3.085 1.715 ;
        RECT  2.855 1.375 3.085 3.240 ;
        RECT  2.855 1.790 5.590 2.020 ;
        RECT  5.250 1.790 5.590 2.220 ;
        RECT  2.855 1.790 3.090 3.240 ;
        RECT  2.750 2.900 3.090 3.240 ;
        RECT  3.860 1.220 4.200 1.560 ;
        RECT  3.860 1.330 6.225 1.560 ;
        RECT  5.940 1.330 6.225 3.140 ;
        RECT  4.470 2.910 6.225 3.140 ;
        RECT  4.470 2.910 4.810 3.250 ;
        RECT  5.120 0.760 5.460 1.100 ;
        RECT  5.120 0.870 6.685 1.100 ;
        RECT  7.375 1.880 8.085 2.220 ;
        RECT  6.455 0.870 6.685 4.180 ;
        RECT  7.375 1.880 7.605 2.940 ;
        RECT  6.455 2.710 7.605 2.940 ;
        RECT  5.010 3.370 6.790 3.600 ;
        RECT  5.010 3.370 5.350 3.995 ;
        RECT  6.455 2.710 6.790 4.180 ;
        RECT  6.450 3.370 6.790 4.180 ;
        RECT  6.915 0.885 9.745 1.115 ;
        RECT  9.515 1.240 10.600 1.580 ;
        RECT  6.915 0.885 7.145 2.480 ;
        RECT  9.515 0.885 9.745 2.920 ;
        RECT  9.670 2.640 10.010 3.470 ;
        RECT  0.115 3.470 3.60 3.700 ;
        RECT  2.855 1.790 4.40 2.020 ;
        RECT  3.860 1.330 5.90 1.560 ;
        RECT  6.915 0.885 8.40 1.115 ;
    END
END NO6I3X4

MACRO NO6I3X2
    CLASS CORE ;
    FOREIGN NO6I3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 2.250 2.395 2.785 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.936  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.580 3.460 8.075 3.850 ;
        RECT  7.580 2.685 7.950 3.850 ;
        RECT  7.720 1.405 7.950 3.850 ;
        RECT  7.390 1.405 7.950 1.690 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.605 1.640 3.655 2.020 ;
        RECT  2.620 1.640 2.905 2.195 ;
        RECT  2.605 1.640 2.905 2.155 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.705 3.560 2.935 ;
        RECT  3.250 2.285 3.560 2.935 ;
        RECT  2.645 2.705 3.025 3.240 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.640 2.060 9.325 2.630 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.120 1.270 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.555 1.625 9.965 2.225 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.360 3.320 8.700 5.280 ;
        RECT  6.800 3.960 7.140 5.280 ;
        RECT  5.520 3.100 5.860 5.280 ;
        RECT  3.715 3.625 4.055 5.280 ;
        RECT  2.300 3.755 2.640 5.280 ;
        RECT  1.290 3.795 1.630 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  9.385 -0.400 9.730 1.040 ;
        RECT  7.990 -0.400 8.330 0.710 ;
        RECT  6.760 -0.400 7.100 0.710 ;
        RECT  3.640 -0.400 3.980 0.950 ;
        RECT  1.380 -0.400 1.720 0.725 ;
        RECT  0.180 -0.400 0.485 0.725 ;
        RECT  0.180 -0.400 0.465 0.755 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.290 1.415 1.135 1.700 ;
        RECT  0.290 1.415 0.520 4.170 ;
        RECT  0.180 3.660 0.520 4.170 ;
        RECT  0.180 3.830 1.060 4.170 ;
        RECT  0.685 0.840 0.970 1.185 ;
        RECT  0.665 0.870 0.970 1.185 ;
        RECT  2.080 0.710 2.420 1.185 ;
        RECT  0.665 0.955 2.420 1.185 ;
        RECT  1.500 0.955 1.730 3.355 ;
        RECT  1.500 3.015 2.140 3.355 ;
        RECT  2.810 0.630 3.150 1.410 ;
        RECT  2.810 1.180 4.115 1.410 ;
        RECT  3.885 1.180 4.115 2.615 ;
        RECT  3.885 2.275 4.360 2.615 ;
        RECT  3.790 2.385 4.020 3.395 ;
        RECT  3.255 3.165 4.020 3.395 ;
        RECT  3.255 3.165 3.485 3.965 ;
        RECT  3.000 3.625 3.485 3.965 ;
        RECT  4.440 1.335 4.830 1.675 ;
        RECT  4.600 1.880 5.620 2.220 ;
        RECT  4.600 1.335 4.830 3.185 ;
        RECT  4.260 2.845 4.830 3.185 ;
        RECT  5.140 0.820 5.480 1.650 ;
        RECT  5.140 1.420 6.080 1.650 ;
        RECT  7.120 2.120 7.490 2.460 ;
        RECT  5.850 1.420 6.080 2.870 ;
        RECT  7.120 2.120 7.350 2.870 ;
        RECT  5.060 2.640 7.350 2.870 ;
        RECT  6.240 2.640 6.580 3.555 ;
        RECT  5.060 2.640 5.290 3.920 ;
        RECT  4.760 3.580 5.290 3.920 ;
        RECT  6.590 0.945 8.410 1.175 ;
        RECT  8.180 1.350 9.130 1.690 ;
        RECT  6.590 0.945 6.820 2.235 ;
        RECT  6.480 1.895 6.820 2.235 ;
        RECT  8.180 0.945 8.410 3.090 ;
        RECT  8.180 2.860 9.890 3.090 ;
        RECT  9.550 2.860 9.890 3.200 ;
        RECT  5.060 2.640 6.60 2.870 ;
    END
END NO6I3X2

MACRO NO6I3X1
    CLASS CORE ;
    FOREIGN NO6I3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.320 3.520 1.810 4.020 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.672  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 3.470 7.435 3.930 ;
        RECT  7.100 1.605 7.330 3.930 ;
        RECT  6.965 1.605 7.330 1.890 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 1.740 2.685 2.070 ;
        RECT  2.015 1.635 2.400 2.025 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.300 3.320 2.630 ;
        RECT  2.960 2.165 3.320 2.630 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.820 1.065 9.325 1.410 ;
        RECT  8.640 1.380 9.055 1.720 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.005 1.290 2.345 ;
        RECT  0.755 2.005 1.090 2.640 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.025 2.250 8.695 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.720 3.885 9.060 5.280 ;
        RECT  6.305 3.035 6.685 5.280 ;
        RECT  4.860 3.615 5.200 5.280 ;
        RECT  3.460 3.910 3.800 5.280 ;
        RECT  2.040 3.060 2.380 5.280 ;
        RECT  1.320 3.060 2.380 3.290 ;
        RECT  1.320 2.720 1.605 3.290 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.925 -0.400 9.270 0.835 ;
        RECT  7.330 -0.400 7.670 0.915 ;
        RECT  6.435 -0.400 6.775 0.880 ;
        RECT  3.680 -0.400 4.020 0.710 ;
        RECT  1.385 -0.400 1.725 0.710 ;
        RECT  0.180 -0.400 0.520 0.690 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.410 1.125 1.695 ;
        RECT  0.180 1.410 0.520 4.200 ;
        RECT  0.180 3.860 1.040 4.200 ;
        RECT  0.635 0.890 0.975 1.180 ;
        RECT  2.085 0.630 2.425 1.180 ;
        RECT  0.635 0.950 2.425 1.180 ;
        RECT  1.555 0.950 1.785 2.490 ;
        RECT  1.555 2.260 2.080 2.490 ;
        RECT  1.850 2.260 2.080 2.830 ;
        RECT  1.850 2.545 2.365 2.830 ;
        RECT  2.690 1.185 3.780 1.510 ;
        RECT  3.550 1.870 4.370 2.210 ;
        RECT  3.550 1.185 3.780 3.140 ;
        RECT  2.760 2.910 3.780 3.140 ;
        RECT  2.760 2.910 3.100 3.880 ;
        RECT  4.020 2.640 4.920 2.925 ;
        RECT  4.480 0.745 5.345 1.090 ;
        RECT  4.805 1.470 5.145 1.930 ;
        RECT  4.805 1.700 5.870 1.930 ;
        RECT  5.635 1.700 5.870 3.875 ;
        RECT  6.585 2.140 6.870 2.480 ;
        RECT  5.635 2.250 6.870 2.480 ;
        RECT  4.100 3.155 5.920 3.385 ;
        RECT  4.100 3.155 4.440 3.760 ;
        RECT  5.635 2.250 5.920 3.875 ;
        RECT  5.580 3.155 5.920 3.875 ;
        RECT  8.130 0.720 8.470 1.060 ;
        RECT  5.865 0.630 6.205 1.375 ;
        RECT  8.130 0.720 8.360 1.375 ;
        RECT  5.865 1.145 8.360 1.375 ;
        RECT  7.565 1.145 7.795 3.275 ;
        RECT  7.565 2.935 8.070 3.275 ;
        RECT  5.865 1.145 7.50 1.375 ;
    END
END NO6I3X1

MACRO NO6I3X0
    CLASS CORE ;
    FOREIGN NO6I3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.040 2.270 2.520 2.685 ;
        RECT  2.040 2.210 2.345 2.685 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.695 1.030 1.135 1.410 ;
        RECT  0.695 0.630 0.925 1.410 ;
        RECT  0.460 0.630 0.925 0.915 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.434  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.860 7.420 3.240 ;
        RECT  7.020 2.710 7.420 3.240 ;
        RECT  7.020 1.475 7.250 3.240 ;
        RECT  6.900 1.475 7.250 1.760 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 2.240 3.605 2.670 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.575 1.480 3.025 2.035 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.650 2.245 8.100 2.790 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.220 0.950 8.695 1.435 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.480 3.530 7.410 5.280 ;
        RECT  5.135 3.610 5.420 5.280 ;
        RECT  3.580 3.500 3.920 5.280 ;
        RECT  2.180 3.520 2.520 5.280 ;
        RECT  0.980 3.410 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.300 -0.400 8.640 0.710 ;
        RECT  6.230 -0.400 7.040 0.715 ;
        RECT  4.140 -0.400 4.480 0.710 ;
        RECT  2.510 -0.400 2.850 0.960 ;
        RECT  1.155 -0.400 1.495 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.160 0.465 3.660 ;
        RECT  0.180 2.100 1.350 2.425 ;
        RECT  0.180 2.100 0.520 3.660 ;
        RECT  1.580 1.160 1.920 1.500 ;
        RECT  1.070 2.725 1.810 3.050 ;
        RECT  1.580 1.160 1.810 3.975 ;
        RECT  1.580 3.635 1.950 3.975 ;
        RECT  3.340 0.630 3.910 0.960 ;
        RECT  3.680 0.630 3.910 1.920 ;
        RECT  3.835 1.690 4.205 2.030 ;
        RECT  3.835 1.690 4.065 3.200 ;
        RECT  2.880 2.970 4.065 3.200 ;
        RECT  2.880 2.970 3.220 3.750 ;
        RECT  4.140 1.170 4.480 1.460 ;
        RECT  4.435 2.160 5.070 2.445 ;
        RECT  4.435 1.225 4.665 2.785 ;
        RECT  4.295 2.590 4.565 2.975 ;
        RECT  4.845 0.745 5.180 1.080 ;
        RECT  4.895 0.745 5.180 1.930 ;
        RECT  4.895 1.700 5.965 1.930 ;
        RECT  5.680 1.700 5.965 3.380 ;
        RECT  5.680 1.990 6.790 2.330 ;
        RECT  4.715 3.150 6.020 3.380 ;
        RECT  5.680 1.990 6.020 3.380 ;
        RECT  4.675 3.185 4.905 3.750 ;
        RECT  4.280 3.410 4.905 3.750 ;
        RECT  5.660 0.630 6.000 1.175 ;
        RECT  7.500 0.630 7.840 1.175 ;
        RECT  5.660 0.945 7.840 1.175 ;
        RECT  7.610 0.630 7.840 1.895 ;
        RECT  7.610 1.665 8.640 1.895 ;
        RECT  8.355 1.665 8.640 3.780 ;
        RECT  8.300 3.440 8.640 3.780 ;
        RECT  5.660 0.945 6.30 1.175 ;
    END
END NO6I3X0

MACRO NO6I2X4
    CLASS CORE ;
    FOREIGN NO6I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.084  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.500 3.825 8.840 4.165 ;
        RECT  8.500 3.540 8.775 4.165 ;
        RECT  7.685 1.345 8.655 1.685 ;
        RECT  7.180 3.540 8.775 3.770 ;
        RECT  7.180 3.430 8.065 3.770 ;
        RECT  7.835 1.345 8.065 3.770 ;
        RECT  7.205 2.660 8.065 3.000 ;
        RECT  7.685 1.345 8.065 3.000 ;
        RECT  7.050 1.345 8.655 1.650 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.310 0.525 3.240 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.210 1.310 2.650 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.185 2.120 10.585 3.240 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.610 1.880 9.955 2.640 ;
        RECT  9.345 1.880 9.955 2.220 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.600 2.250 4.285 2.650 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.685 2.250 3.270 2.750 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 3.470 10.530 5.280 ;
        RECT  7.740 4.170 8.080 5.280 ;
        RECT  6.620 4.170 6.960 5.280 ;
        RECT  5.100 3.830 5.440 5.280 ;
        RECT  2.690 3.610 3.030 5.280 ;
        RECT  1.300 3.650 1.640 5.280 ;
        RECT  0.180 3.650 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 0.715 ;
        RECT  9.070 -0.400 9.410 0.655 ;
        RECT  7.810 -0.400 8.150 0.655 ;
        RECT  6.290 -0.400 6.630 0.655 ;
        RECT  3.790 -0.400 4.130 0.720 ;
        RECT  2.650 -0.400 2.990 0.720 ;
        RECT  1.190 -0.400 1.530 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.360 0.520 1.700 ;
        RECT  0.180 1.470 1.770 1.700 ;
        RECT  1.540 2.260 1.995 2.600 ;
        RECT  1.540 1.470 1.770 3.220 ;
        RECT  0.755 2.880 1.770 3.220 ;
        RECT  2.000 1.235 2.455 1.575 ;
        RECT  2.225 1.790 4.960 2.020 ;
        RECT  4.620 1.790 4.960 2.220 ;
        RECT  2.225 1.235 2.455 3.335 ;
        RECT  2.060 2.995 2.455 3.335 ;
        RECT  3.230 1.220 3.570 1.560 ;
        RECT  3.230 1.330 5.595 1.560 ;
        RECT  5.310 1.330 5.595 3.140 ;
        RECT  3.840 2.910 5.595 3.140 ;
        RECT  3.840 2.910 4.180 3.305 ;
        RECT  4.490 0.760 4.830 1.100 ;
        RECT  4.490 0.870 6.055 1.100 ;
        RECT  6.745 1.880 7.455 2.220 ;
        RECT  5.825 0.870 6.055 4.180 ;
        RECT  6.745 1.880 6.975 2.950 ;
        RECT  5.825 2.710 6.975 2.950 ;
        RECT  4.490 3.370 6.160 3.600 ;
        RECT  4.490 3.370 4.720 3.995 ;
        RECT  4.380 3.655 4.720 3.995 ;
        RECT  5.825 2.710 6.160 4.180 ;
        RECT  5.820 3.370 6.160 4.180 ;
        RECT  6.285 0.885 9.115 1.115 ;
        RECT  8.885 1.240 9.970 1.580 ;
        RECT  6.285 0.885 6.515 2.480 ;
        RECT  8.885 0.885 9.115 2.920 ;
        RECT  9.040 2.640 9.380 3.470 ;
        RECT  2.225 1.790 3.40 2.020 ;
        RECT  3.230 1.330 4.60 1.560 ;
        RECT  6.285 0.885 8.50 1.115 ;
    END
END NO6I2X4

MACRO NO6I2X2
    CLASS CORE ;
    FOREIGN NO6I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.936  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 3.460 7.445 3.850 ;
        RECT  6.950 2.685 7.320 3.850 ;
        RECT  7.090 1.405 7.320 3.850 ;
        RECT  6.760 1.405 7.320 1.690 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.640 3.025 2.020 ;
        RECT  1.990 1.640 2.275 2.195 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.705 2.930 2.935 ;
        RECT  2.620 2.285 2.930 2.935 ;
        RECT  2.015 2.705 2.395 3.240 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.010 2.060 8.695 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.600 0.550 2.220 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.240 2.250 1.765 2.690 ;
        RECT  1.240 2.120 1.760 2.690 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.925 1.625 9.335 2.225 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.730 3.320 8.070 5.280 ;
        RECT  6.170 4.080 6.510 5.280 ;
        RECT  4.890 3.100 5.230 5.280 ;
        RECT  3.085 3.660 3.425 5.280 ;
        RECT  1.445 2.920 1.785 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.755 -0.400 9.100 1.040 ;
        RECT  7.360 -0.400 7.700 0.710 ;
        RECT  6.130 -0.400 6.470 0.710 ;
        RECT  3.010 -0.400 3.350 0.950 ;
        RECT  1.380 -0.400 1.720 1.050 ;
        RECT  0.180 -0.400 0.520 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.360 1.135 1.700 ;
        RECT  0.180 2.775 1.010 3.115 ;
        RECT  0.780 1.360 1.010 4.170 ;
        RECT  0.780 3.830 1.125 4.170 ;
        RECT  2.180 0.630 2.520 1.410 ;
        RECT  2.180 1.180 3.485 1.410 ;
        RECT  3.255 1.180 3.485 2.615 ;
        RECT  3.255 2.275 3.730 2.615 ;
        RECT  3.160 2.385 3.390 3.430 ;
        RECT  2.625 3.200 3.390 3.430 ;
        RECT  2.625 3.200 2.855 4.000 ;
        RECT  2.370 3.660 2.855 4.000 ;
        RECT  3.810 1.335 4.200 1.675 ;
        RECT  3.970 1.880 4.990 2.220 ;
        RECT  3.970 1.335 4.200 3.220 ;
        RECT  3.630 2.880 4.200 3.220 ;
        RECT  4.510 0.820 4.850 1.650 ;
        RECT  4.510 1.420 5.450 1.650 ;
        RECT  6.490 2.120 6.860 2.460 ;
        RECT  5.220 1.420 5.450 2.870 ;
        RECT  6.490 2.120 6.720 2.870 ;
        RECT  4.430 2.640 6.720 2.870 ;
        RECT  5.610 2.640 5.950 3.555 ;
        RECT  4.430 2.640 4.660 3.960 ;
        RECT  4.130 3.620 4.660 3.960 ;
        RECT  5.960 0.945 7.780 1.175 ;
        RECT  7.550 1.350 8.500 1.690 ;
        RECT  5.960 0.945 6.190 2.235 ;
        RECT  5.850 1.895 6.190 2.235 ;
        RECT  7.550 0.945 7.780 3.090 ;
        RECT  7.550 2.860 9.260 3.090 ;
        RECT  8.920 2.860 9.260 3.200 ;
        RECT  4.430 2.640 5.20 2.870 ;
    END
END NO6I2X2

MACRO NO6I2X1
    CLASS CORE ;
    FOREIGN NO6I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.672  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.420 3.470 6.805 3.930 ;
        RECT  6.485 1.605 6.715 3.930 ;
        RECT  6.375 1.605 6.715 1.890 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.740 2.095 2.065 ;
        RECT  1.385 1.640 1.765 2.065 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.295 2.670 2.655 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.900 0.970 1.150 ;
        RECT  0.660 0.840 0.970 1.150 ;
        RECT  0.630 0.860 0.970 1.150 ;
        RECT  0.125 0.900 0.505 1.410 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.020 1.640 8.695 2.020 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.305 1.445 2.645 ;
        RECT  0.755 2.305 1.115 3.240 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.405 2.250 8.065 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.260 2.975 8.600 5.280 ;
        RECT  5.675 3.035 6.055 5.280 ;
        RECT  4.230 3.615 4.570 5.280 ;
        RECT  2.630 3.645 2.970 5.280 ;
        RECT  1.345 2.890 1.685 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.295 -0.400 8.640 1.055 ;
        RECT  6.700 -0.400 7.040 0.915 ;
        RECT  5.825 -0.400 6.165 0.880 ;
        RECT  3.070 -0.400 3.410 0.710 ;
        RECT  1.380 -0.400 1.720 0.925 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        RECT  0.180 -0.400 0.500 0.670 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.380 1.120 1.890 ;
        RECT  0.180 1.660 1.120 1.890 ;
        RECT  0.180 1.660 0.520 4.250 ;
        RECT  2.080 1.185 3.150 1.510 ;
        RECT  2.920 1.750 3.765 2.090 ;
        RECT  2.920 1.185 3.150 3.245 ;
        RECT  2.065 2.905 3.150 3.245 ;
        RECT  3.390 2.640 4.290 2.925 ;
        RECT  3.870 0.745 4.735 1.090 ;
        RECT  4.195 1.470 4.535 1.930 ;
        RECT  4.195 1.700 5.240 1.930 ;
        RECT  5.005 1.700 5.240 3.875 ;
        RECT  5.005 2.140 6.255 2.480 ;
        RECT  3.470 3.155 5.290 3.385 ;
        RECT  3.470 3.155 3.810 3.760 ;
        RECT  5.005 2.140 5.290 3.875 ;
        RECT  4.950 3.155 5.290 3.875 ;
        RECT  5.255 0.630 5.595 1.375 ;
        RECT  7.500 0.720 7.840 1.375 ;
        RECT  5.255 1.145 7.840 1.375 ;
        RECT  6.945 1.145 7.175 3.275 ;
        RECT  6.945 2.935 7.450 3.275 ;
        RECT  5.255 1.145 6.60 1.375 ;
    END
END NO6I2X1

MACRO NO6I2X0
    CLASS CORE ;
    FOREIGN NO6I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.410 2.250 1.765 2.815 ;
        RECT  1.410 2.210 1.730 2.815 ;
        RECT  1.410 2.035 1.715 2.815 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.630 0.720 2.125 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.434  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.860 6.790 3.240 ;
        RECT  6.390 2.710 6.790 3.240 ;
        RECT  6.390 1.405 6.620 3.240 ;
        RECT  6.270 1.405 6.620 1.750 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.440 2.360 2.975 2.670 ;
        RECT  2.620 2.185 2.975 2.670 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 1.545 2.390 2.100 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.020 2.245 7.470 2.790 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.590 0.950 8.065 1.435 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  5.850 3.530 6.780 5.280 ;
        RECT  4.505 3.675 4.790 5.280 ;
        RECT  2.950 3.430 3.290 5.280 ;
        RECT  1.550 3.450 1.890 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 0.710 ;
        RECT  5.600 -0.400 6.410 0.715 ;
        RECT  3.510 -0.400 3.850 0.710 ;
        RECT  1.880 -0.400 2.220 0.960 ;
        RECT  0.345 -0.400 0.690 0.855 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.950 1.160 1.290 1.500 ;
        RECT  0.440 2.640 1.180 2.980 ;
        RECT  0.950 1.160 1.180 3.975 ;
        RECT  0.950 3.635 1.320 3.975 ;
        RECT  2.710 0.630 3.280 0.960 ;
        RECT  3.050 0.630 3.280 1.915 ;
        RECT  3.205 1.690 3.575 2.030 ;
        RECT  3.205 1.690 3.435 3.130 ;
        RECT  2.250 2.900 3.435 3.130 ;
        RECT  2.250 2.900 2.590 3.750 ;
        RECT  3.510 1.170 3.850 1.455 ;
        RECT  3.805 2.160 4.440 2.445 ;
        RECT  3.805 1.225 4.035 2.820 ;
        RECT  3.665 2.520 3.935 3.050 ;
        RECT  4.215 0.745 4.550 1.080 ;
        RECT  4.265 0.745 4.550 1.930 ;
        RECT  4.265 1.700 5.335 1.930 ;
        RECT  5.050 1.700 5.335 3.445 ;
        RECT  5.050 1.990 6.160 2.330 ;
        RECT  4.110 3.215 5.390 3.445 ;
        RECT  5.050 1.990 5.390 3.445 ;
        RECT  4.045 3.275 4.275 3.800 ;
        RECT  3.650 3.460 4.275 3.800 ;
        RECT  5.030 0.630 5.370 1.175 ;
        RECT  6.870 0.630 7.210 1.175 ;
        RECT  5.030 0.945 7.210 1.175 ;
        RECT  5.030 0.945 6.40 1.175 ;
        RECT  6.980 0.630 7.210 1.895 ;
        RECT  6.980 1.665 8.010 1.895 ;
        RECT  7.725 1.665 8.010 3.780 ;
        RECT  7.670 3.440 8.010 3.780 ;
    END
END NO6I2X0

MACRO NO6I1X4
    CLASS CORE ;
    FOREIGN NO6I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.084  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.500 3.825 8.840 4.165 ;
        RECT  8.500 3.540 8.730 4.165 ;
        RECT  7.685 1.345 8.655 1.685 ;
        RECT  7.180 3.540 8.730 3.770 ;
        RECT  7.180 3.430 8.065 3.770 ;
        RECT  7.835 1.345 8.065 3.770 ;
        RECT  7.205 2.660 8.065 3.000 ;
        RECT  7.685 1.345 8.065 3.000 ;
        RECT  7.050 1.345 8.655 1.650 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.440 0.770 3.850 ;
        END
    END AN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.185 2.120 10.585 3.240 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.240 2.860 1.765 3.240 ;
        RECT  1.240 2.310 1.615 3.240 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.610 1.880 9.955 2.650 ;
        RECT  9.345 1.880 9.955 2.220 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.600 2.250 4.285 2.650 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.195 3.655 3.850 ;
        RECT  2.940 3.195 3.655 3.425 ;
        RECT  2.940 2.310 3.270 3.425 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 3.470 10.530 5.280 ;
        RECT  7.740 4.170 8.080 5.280 ;
        RECT  6.620 4.170 6.960 5.280 ;
        RECT  5.100 3.830 5.440 5.280 ;
        RECT  2.690 3.655 3.030 5.280 ;
        RECT  1.000 3.470 1.340 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 0.715 ;
        RECT  9.070 -0.400 9.410 0.655 ;
        RECT  7.810 -0.400 8.150 0.655 ;
        RECT  6.290 -0.400 6.630 0.655 ;
        RECT  3.790 -0.400 4.130 0.720 ;
        RECT  2.450 -0.400 2.790 1.160 ;
        RECT  0.910 -0.400 1.250 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.240 1.360 0.630 2.080 ;
        RECT  0.240 1.850 2.250 2.080 ;
        RECT  1.910 1.850 2.250 2.220 ;
        RECT  0.240 1.360 0.580 3.210 ;
        RECT  1.690 1.280 2.030 1.620 ;
        RECT  1.690 1.390 2.710 1.620 ;
        RECT  2.480 1.790 4.960 2.020 ;
        RECT  4.620 1.790 4.960 2.220 ;
        RECT  2.480 1.390 2.710 3.320 ;
        RECT  2.150 2.980 2.710 3.320 ;
        RECT  3.230 1.220 3.570 1.560 ;
        RECT  3.230 1.330 5.595 1.560 ;
        RECT  5.310 1.330 5.595 3.140 ;
        RECT  3.885 2.910 5.595 3.140 ;
        RECT  3.885 2.910 4.180 3.305 ;
        RECT  4.490 0.760 4.830 1.100 ;
        RECT  4.490 0.870 6.055 1.100 ;
        RECT  6.745 1.880 7.280 2.220 ;
        RECT  5.825 0.870 6.055 4.180 ;
        RECT  6.745 1.880 6.975 2.940 ;
        RECT  5.825 2.710 6.975 2.940 ;
        RECT  4.490 3.370 6.160 3.600 ;
        RECT  4.490 3.370 4.720 3.995 ;
        RECT  4.380 3.655 4.720 3.995 ;
        RECT  5.825 2.710 6.160 4.180 ;
        RECT  5.820 3.370 6.160 4.180 ;
        RECT  6.285 0.885 9.115 1.115 ;
        RECT  8.885 1.240 9.970 1.580 ;
        RECT  6.285 0.885 6.515 2.480 ;
        RECT  8.885 0.885 9.115 2.920 ;
        RECT  9.040 2.640 9.380 3.470 ;
        RECT  0.240 1.850 1.80 2.080 ;
        RECT  2.480 1.790 3.80 2.020 ;
        RECT  3.230 1.330 4.70 1.560 ;
        RECT  6.285 0.885 8.00 1.115 ;
    END
END NO6I1X4

MACRO NO6I1X2
    CLASS CORE ;
    FOREIGN NO6I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.936  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 3.460 7.445 3.850 ;
        RECT  6.950 2.685 7.320 3.850 ;
        RECT  7.090 1.405 7.320 3.850 ;
        RECT  6.760 1.405 7.320 1.690 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.585 2.250 4.285 2.655 ;
        END
    END AN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.060 8.220 2.630 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.690 3.470 2.395 4.055 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.600 0.550 2.195 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.240 1.910 1.765 2.250 ;
        RECT  1.385 1.640 1.765 2.250 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.925 1.625 9.335 2.225 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.730 2.860 8.070 5.280 ;
        RECT  6.170 4.080 6.510 5.280 ;
        RECT  4.940 3.275 5.230 5.280 ;
        RECT  4.945 3.220 5.230 5.280 ;
        RECT  3.630 3.540 3.970 5.280 ;
        RECT  1.120 3.660 1.460 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.755 -0.400 9.100 1.040 ;
        RECT  7.360 -0.400 7.700 0.710 ;
        RECT  6.130 -0.400 6.470 0.710 ;
        RECT  2.780 -0.400 3.120 0.655 ;
        RECT  1.380 -0.400 1.720 1.025 ;
        RECT  0.180 -0.400 0.520 1.025 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.335 1.120 1.675 ;
        RECT  0.780 1.335 1.010 3.070 ;
        RECT  0.180 2.730 1.010 3.070 ;
        RECT  0.545 2.730 0.890 4.170 ;
        RECT  3.400 1.345 3.745 2.020 ;
        RECT  2.455 1.790 3.745 2.020 ;
        RECT  2.455 1.790 3.355 2.195 ;
        RECT  3.125 1.790 3.355 3.960 ;
        RECT  2.870 3.620 3.355 3.960 ;
        RECT  1.995 0.685 2.420 1.115 ;
        RECT  1.995 0.885 4.205 1.115 ;
        RECT  3.975 0.885 4.205 2.020 ;
        RECT  3.975 1.790 4.990 2.020 ;
        RECT  4.650 1.790 4.990 2.220 ;
        RECT  1.995 0.685 2.225 3.100 ;
        RECT  1.995 2.760 2.895 3.100 ;
        RECT  4.510 0.805 4.850 1.560 ;
        RECT  4.510 1.330 5.450 1.560 ;
        RECT  6.490 2.120 6.860 2.460 ;
        RECT  5.220 1.330 5.450 2.980 ;
        RECT  5.220 2.640 6.720 2.870 ;
        RECT  6.490 2.120 6.720 2.870 ;
        RECT  4.505 2.725 5.950 2.980 ;
        RECT  4.130 2.885 4.715 3.225 ;
        RECT  5.610 2.640 5.950 3.555 ;
        RECT  5.960 0.945 8.390 1.175 ;
        RECT  8.160 0.945 8.390 1.690 ;
        RECT  8.160 1.350 8.695 1.690 ;
        RECT  5.960 0.945 6.190 2.235 ;
        RECT  5.850 1.895 6.190 2.235 ;
        RECT  8.465 1.350 8.695 3.110 ;
        RECT  8.465 2.770 9.260 3.110 ;
        RECT  1.995 0.885 3.60 1.115 ;
        RECT  5.960 0.945 7.50 1.175 ;
    END
END NO6I1X2

MACRO NO6I1X1
    CLASS CORE ;
    FOREIGN NO6I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.065 1.680 2.395 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.672  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.420 3.735 6.875 4.075 ;
        RECT  6.420 3.470 6.820 4.075 ;
        RECT  6.555 1.470 6.785 4.075 ;
        RECT  6.445 1.470 6.785 1.790 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.530 1.660 4.295 1.970 ;
        RECT  3.530 1.640 3.875 1.970 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.900 0.970 1.150 ;
        RECT  0.660 0.840 0.970 1.150 ;
        RECT  0.630 0.860 0.970 1.150 ;
        RECT  0.125 0.900 0.505 1.410 ;
        END
    END C
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.150 1.600 8.705 2.025 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.905 2.100 1.375 2.385 ;
        RECT  0.755 2.860 1.135 3.240 ;
        RECT  0.905 2.100 1.135 3.240 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.520 2.245 8.080 2.680 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.270 3.885 8.610 5.280 ;
        RECT  5.815 3.230 6.155 5.280 ;
        RECT  4.330 3.615 4.670 5.280 ;
        RECT  3.090 2.660 3.395 5.280 ;
        RECT  3.055 2.660 3.395 3.585 ;
        RECT  1.365 3.910 1.710 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.295 -0.400 8.640 0.780 ;
        RECT  6.845 -0.400 7.185 0.780 ;
        RECT  5.825 -0.400 6.165 0.780 ;
        RECT  2.780 -0.400 3.120 0.710 ;
        RECT  1.380 -0.400 1.720 0.875 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        RECT  0.180 -0.400 0.500 0.670 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.380 1.120 1.870 ;
        RECT  0.180 1.640 1.120 1.870 ;
        RECT  0.180 1.640 0.520 4.250 ;
        RECT  2.180 1.070 2.530 1.410 ;
        RECT  1.605 1.120 2.530 1.410 ;
        RECT  1.605 1.120 1.835 3.310 ;
        RECT  1.605 3.080 2.740 3.310 ;
        RECT  2.400 3.080 2.740 4.100 ;
        RECT  2.400 3.760 2.860 4.100 ;
        RECT  3.580 0.630 3.920 0.950 ;
        RECT  3.580 0.630 3.820 1.335 ;
        RECT  3.070 1.105 3.820 1.335 ;
        RECT  3.070 1.105 3.300 2.430 ;
        RECT  2.700 1.965 3.300 2.305 ;
        RECT  3.070 2.200 4.115 2.430 ;
        RECT  3.775 2.200 4.115 2.900 ;
        RECT  4.195 1.145 5.305 1.430 ;
        RECT  5.070 1.145 5.305 3.875 ;
        RECT  5.965 2.660 6.305 3.000 ;
        RECT  5.070 2.770 6.305 3.000 ;
        RECT  3.625 3.155 5.390 3.385 ;
        RECT  3.625 3.155 3.910 3.760 ;
        RECT  5.070 2.770 5.390 3.875 ;
        RECT  5.050 3.155 5.390 3.875 ;
        RECT  5.645 1.010 7.985 1.240 ;
        RECT  7.060 1.010 7.985 1.430 ;
        RECT  5.645 1.010 5.875 2.325 ;
        RECT  5.535 1.985 5.875 2.325 ;
        RECT  7.060 1.010 7.290 3.275 ;
        RECT  7.060 2.935 7.620 3.275 ;
        RECT  5.645 1.010 6.60 1.240 ;
    END
END NO6I1X1

MACRO NO6I1X0
    CLASS CORE ;
    FOREIGN NO6I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.640 2.050 1.135 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.040 1.115 ;
        RECT  0.750 0.630 1.040 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.860 6.790 3.240 ;
        RECT  6.390 2.710 6.790 3.240 ;
        RECT  6.390 1.485 6.620 3.240 ;
        RECT  6.270 1.485 6.620 1.770 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.955 1.845 3.385 2.185 ;
        RECT  2.645 1.640 3.150 2.020 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 2.025 1.750 2.660 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.020 2.200 7.425 2.750 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.590 0.950 8.065 1.435 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  5.850 3.530 6.780 5.280 ;
        RECT  4.510 3.580 4.795 5.280 ;
        RECT  2.915 3.360 3.255 5.280 ;
        RECT  1.270 3.485 1.610 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 0.710 ;
        RECT  5.600 -0.400 6.410 0.715 ;
        RECT  2.780 -0.400 3.120 0.690 ;
        RECT  1.380 -0.400 1.720 0.960 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.630 ;
        RECT  0.180 1.590 0.965 1.820 ;
        RECT  0.180 1.590 0.410 3.825 ;
        RECT  0.180 3.485 0.930 3.825 ;
        RECT  0.700 3.635 1.040 3.975 ;
        RECT  3.380 1.380 3.845 1.615 ;
        RECT  2.440 2.285 2.725 2.645 ;
        RECT  2.440 2.415 3.845 2.645 ;
        RECT  3.615 1.380 3.845 2.970 ;
        RECT  3.515 2.415 3.845 2.970 ;
        RECT  1.980 0.630 2.420 1.150 ;
        RECT  3.660 0.805 4.000 1.150 ;
        RECT  1.980 0.920 4.000 1.150 ;
        RECT  1.980 0.630 2.210 3.825 ;
        RECT  1.980 3.485 2.555 3.825 ;
        RECT  4.230 0.745 4.550 1.635 ;
        RECT  4.230 1.405 5.335 1.635 ;
        RECT  5.050 1.405 5.335 3.280 ;
        RECT  5.050 1.990 6.160 2.330 ;
        RECT  4.100 3.050 5.390 3.280 ;
        RECT  5.050 1.990 5.390 3.280 ;
        RECT  4.050 3.085 4.280 3.680 ;
        RECT  3.650 3.340 4.280 3.680 ;
        RECT  5.030 0.630 5.370 1.175 ;
        RECT  6.870 0.665 7.210 1.175 ;
        RECT  5.030 0.945 7.210 1.175 ;
        RECT  6.980 0.665 7.210 1.950 ;
        RECT  6.980 1.720 8.010 1.950 ;
        RECT  7.670 1.720 8.010 3.780 ;
        RECT  1.980 0.920 3.60 1.150 ;
        RECT  5.030 0.945 6.30 1.175 ;
    END
END NO6I1X0

MACRO NO5X4
    CLASS CORE ;
    FOREIGN NO5X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 1.040 8.015 4.160 ;
        RECT  6.470 2.205 8.015 2.655 ;
        RECT  6.230 3.115 6.700 4.160 ;
        RECT  6.470 1.040 6.700 4.160 ;
        RECT  6.230 1.040 6.700 1.380 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 3.025 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.910 3.890 4.250 ;
        RECT  3.275 3.470 3.655 4.250 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.860 1.135 3.240 ;
        RECT  0.750 2.135 0.980 3.240 ;
        RECT  0.575 2.135 0.980 2.480 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.910 1.530 2.395 2.020 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 2.250 1.765 2.625 ;
        RECT  1.210 1.780 1.520 2.625 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.950 -0.400 7.290 1.510 ;
        RECT  5.470 -0.400 5.810 1.000 ;
        RECT  3.620 -0.400 3.960 0.710 ;
        RECT  2.380 -0.400 2.720 0.710 ;
        RECT  0.900 -0.400 1.240 1.040 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.950 2.920 7.290 5.280 ;
        RECT  5.510 3.180 5.850 5.280 ;
        RECT  4.120 2.720 4.370 5.280 ;
        RECT  4.030 2.720 4.370 3.600 ;
        RECT  1.960 2.860 2.290 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.970 1.400 3.620 1.715 ;
        RECT  3.270 2.150 4.865 2.490 ;
        RECT  3.270 1.400 3.620 3.240 ;
        RECT  1.470 0.940 4.090 1.170 ;
        RECT  0.115 0.735 0.520 1.500 ;
        RECT  1.470 0.940 1.960 1.280 ;
        RECT  0.115 1.270 1.700 1.430 ;
        RECT  0.115 1.270 1.675 1.500 ;
        RECT  3.860 0.940 4.090 1.920 ;
        RECT  3.860 1.690 5.460 1.920 ;
        RECT  5.230 1.690 5.460 2.490 ;
        RECT  5.230 2.150 5.565 2.490 ;
        RECT  0.115 0.735 0.345 4.175 ;
        RECT  0.115 2.715 0.520 4.175 ;
        RECT  4.320 0.700 4.660 1.460 ;
        RECT  4.320 1.230 6.000 1.460 ;
        RECT  5.770 1.230 6.000 2.040 ;
        RECT  5.795 1.890 6.240 2.230 ;
        RECT  5.795 1.890 6.060 2.950 ;
        RECT  4.750 2.720 6.060 2.950 ;
        RECT  4.750 2.720 5.090 4.180 ;
        RECT  1.470 0.940 3.20 1.170 ;
    END
END NO5X4

MACRO NO5X2
    CLASS CORE ;
    FOREIGN NO5X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.280  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.675 2.040 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.315 2.320 1.715 3.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.590 2.225 1.085 2.685 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.280  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.785 2.250 6.355 2.705 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.375 2.250 4.925 2.630 ;
        RECT  4.330 3.040 4.670 3.960 ;
        RECT  4.375 2.250 4.670 3.960 ;
        RECT  4.375 1.680 4.605 3.960 ;
        RECT  4.230 1.680 4.605 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.306  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 2.240 2.395 2.750 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.105 2.985 5.445 5.280 ;
        RECT  3.610 3.080 3.950 5.280 ;
        RECT  2.170 3.040 2.510 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 0.950 ;
        RECT  4.890 -0.400 5.230 0.950 ;
        RECT  2.340 -0.400 2.680 1.430 ;
        RECT  0.900 -0.400 1.240 1.430 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.180 0.520 1.945 ;
        RECT  1.620 1.180 1.960 1.945 ;
        RECT  0.115 1.715 2.900 1.945 ;
        RECT  2.575 1.715 2.900 2.060 ;
        RECT  0.115 1.180 0.360 3.240 ;
        RECT  0.350 2.990 0.690 3.955 ;
        RECT  3.130 0.700 3.870 0.990 ;
        RECT  3.130 0.700 3.360 2.850 ;
        RECT  2.890 2.520 4.145 2.850 ;
        RECT  2.890 2.520 3.230 3.960 ;
        RECT  5.650 1.060 5.990 1.410 ;
        RECT  4.745 1.180 6.815 1.410 ;
        RECT  3.590 1.220 4.935 1.450 ;
        RECT  3.590 1.220 3.930 2.070 ;
        RECT  6.585 1.180 6.815 3.255 ;
        RECT  6.255 3.000 6.595 3.960 ;
        RECT  0.115 1.715 1.40 1.945 ;
        RECT  4.745 1.180 5.80 1.410 ;
    END
END NO5X2

MACRO NO5X1
    CLASS CORE ;
    FOREIGN NO5X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.660 2.120 1.135 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.730 2.025 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.890 2.435 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 1.690 1.765 3.240 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.250 6.355 2.630 ;
        RECT  6.070 2.025 6.355 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.815 1.030 3.655 1.420 ;
        RECT  2.960 2.640 3.300 3.560 ;
        RECT  2.815 1.030 3.045 2.870 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.160 2.670 5.500 5.280 ;
        RECT  3.680 2.640 4.020 5.280 ;
        RECT  2.240 2.885 2.585 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.100 -0.400 6.640 0.710 ;
        RECT  0.980 -0.400 2.595 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.120 1.995 1.460 ;
        RECT  0.180 1.120 0.410 3.205 ;
        RECT  0.180 2.920 1.005 3.205 ;
        RECT  0.470 2.920 1.005 3.260 ;
        RECT  0.470 2.920 0.810 3.965 ;
        RECT  3.910 1.095 4.250 2.055 ;
        RECT  3.275 1.715 4.250 2.055 ;
        RECT  3.275 1.770 4.780 2.055 ;
        RECT  4.440 1.770 4.780 3.015 ;
        RECT  4.150 0.630 4.835 0.865 ;
        RECT  4.605 0.630 4.835 1.410 ;
        RECT  4.605 1.070 6.815 1.410 ;
        RECT  6.585 1.070 6.815 3.200 ;
        RECT  6.310 2.860 6.815 3.200 ;
        RECT  6.310 2.860 6.540 4.150 ;
        RECT  5.890 3.810 6.540 4.150 ;
        RECT  4.605 1.070 5.40 1.410 ;
    END
END NO5X1

MACRO NO5X0
    CLASS CORE ;
    FOREIGN NO5X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.660 2.240 1.135 2.755 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.740 5.725 2.080 ;
        RECT  4.535 1.640 4.915 2.080 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.300 6.355 2.630 ;
        RECT  6.070 2.160 6.355 2.630 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.115 2.435 2.695 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 1.840 1.765 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.800 1.030 3.655 1.460 ;
        RECT  2.980 2.390 3.320 3.360 ;
        RECT  2.800 1.030 3.030 2.705 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.380 3.670 5.720 5.280 ;
        RECT  3.780 3.020 4.120 5.280 ;
        RECT  2.280 3.040 2.625 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.100 -0.400 6.640 0.710 ;
        RECT  0.980 -0.400 2.595 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.120 1.995 1.460 ;
        RECT  0.180 1.120 0.410 3.325 ;
        RECT  0.180 3.040 0.965 3.325 ;
        RECT  0.470 3.040 0.965 3.380 ;
        RECT  0.470 3.040 0.810 3.940 ;
        RECT  3.885 1.175 4.210 2.055 ;
        RECT  3.260 1.715 4.210 2.055 ;
        RECT  3.925 1.175 4.210 2.690 ;
        RECT  3.925 2.460 4.920 2.690 ;
        RECT  4.580 2.460 4.920 3.360 ;
        RECT  4.150 0.630 4.825 0.945 ;
        RECT  4.595 0.630 4.825 1.300 ;
        RECT  4.595 1.070 6.815 1.300 ;
        RECT  5.685 1.070 6.815 1.410 ;
        RECT  6.585 1.070 6.815 3.360 ;
        RECT  6.410 3.020 6.640 4.250 ;
        RECT  5.950 3.910 6.640 4.250 ;
        RECT  4.595 1.070 5.90 1.300 ;
    END
END NO5X0

MACRO NO5I4X4
    CLASS CORE ;
    FOREIGN NO5I4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.660 3.450 2.395 3.850 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.940 3.235 9.325 3.850 ;
        RECT  8.740 3.235 9.325 3.575 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.480 3.370 6.980 4.180 ;
        RECT  6.480 2.660 6.710 4.180 ;
        RECT  4.990 1.345 6.650 1.630 ;
        RECT  5.320 2.660 6.710 2.890 ;
        RECT  5.795 1.345 6.175 2.890 ;
        RECT  5.320 2.660 5.660 3.770 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.065 0.525 2.740 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.880 1.315 2.220 ;
        RECT  0.755 1.880 1.135 2.630 ;
        END
    END BN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.140 1.030 8.695 1.410 ;
        RECT  8.140 0.630 8.370 1.410 ;
        RECT  7.810 0.630 8.370 0.940 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.370 3.805 8.710 5.280 ;
        RECT  5.880 4.170 6.220 5.280 ;
        RECT  4.760 4.170 5.100 5.280 ;
        RECT  3.280 3.655 3.620 5.280 ;
        RECT  1.980 4.080 2.320 5.280 ;
        RECT  0.880 3.650 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.600 -0.400 8.945 0.800 ;
        RECT  7.010 -0.400 7.350 0.655 ;
        RECT  5.750 -0.400 6.090 0.655 ;
        RECT  4.230 -0.400 4.570 0.655 ;
        RECT  1.525 -0.400 1.865 0.960 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.095 0.630 2.600 0.940 ;
        RECT  0.225 0.630 0.565 1.440 ;
        RECT  2.095 0.630 2.325 1.440 ;
        RECT  0.225 1.210 2.325 1.440 ;
        RECT  1.420 2.880 1.775 3.220 ;
        RECT  1.545 1.210 1.775 3.220 ;
        RECT  0.290 2.990 1.775 3.220 ;
        RECT  0.290 2.990 0.520 4.155 ;
        RECT  0.180 3.815 0.520 4.155 ;
        RECT  2.555 1.345 3.080 1.685 ;
        RECT  2.740 2.140 3.500 2.480 ;
        RECT  2.740 1.345 3.080 3.170 ;
        RECT  3.040 0.700 3.380 1.040 ;
        RECT  3.040 0.810 3.960 1.040 ;
        RECT  4.860 1.860 5.565 2.200 ;
        RECT  3.730 0.810 3.960 2.940 ;
        RECT  4.860 1.860 5.090 2.940 ;
        RECT  3.730 2.710 5.090 2.940 ;
        RECT  4.000 2.710 4.340 4.180 ;
        RECT  4.300 0.885 7.190 1.115 ;
        RECT  6.960 1.240 7.910 1.580 ;
        RECT  4.300 0.885 4.530 2.480 ;
        RECT  4.190 2.140 4.530 2.480 ;
        RECT  6.960 0.885 7.190 3.020 ;
        RECT  6.960 2.690 7.520 3.020 ;
        RECT  7.420 2.120 9.270 2.350 ;
        RECT  7.420 2.120 7.760 2.460 ;
        RECT  8.930 1.340 9.270 3.005 ;
        RECT  0.225 1.210 1.50 1.440 ;
        RECT  4.300 0.885 6.60 1.115 ;
    END
END NO5I4X4

MACRO NO5I4X2
    CLASS CORE ;
    FOREIGN NO5I4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.955 1.590 4.425 2.110 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.850 7.500 3.765 ;
        RECT  7.270 1.240 7.500 3.765 ;
        RECT  7.110 1.240 7.500 1.580 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 1.745 2.690 2.070 ;
        RECT  2.035 1.630 2.405 2.030 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.300 3.265 2.640 ;
        RECT  2.950 2.190 3.265 2.640 ;
        END
    END BN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.320 3.520 1.810 4.020 ;
        END
    END DN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.005 1.290 2.345 ;
        RECT  0.755 2.005 1.135 2.580 ;
        RECT  0.755 2.005 1.110 2.605 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.670 4.170 8.010 5.280 ;
        RECT  6.390 2.960 6.730 5.280 ;
        RECT  4.950 3.590 5.290 5.280 ;
        RECT  3.460 3.380 3.800 5.280 ;
        RECT  2.040 3.060 2.380 5.280 ;
        RECT  1.290 3.060 2.380 3.290 ;
        RECT  1.290 2.750 1.605 3.290 ;
        RECT  1.320 2.720 1.605 3.290 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 0.720 ;
        RECT  6.550 -0.400 6.890 0.720 ;
        RECT  4.100 -0.400 4.440 0.710 ;
        RECT  1.380 -0.400 1.720 0.710 ;
        RECT  0.180 -0.400 0.520 0.670 ;
        RECT  0.180 -0.400 0.495 0.690 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.410 1.120 1.695 ;
        RECT  0.180 1.410 0.520 4.200 ;
        RECT  0.180 3.860 1.040 4.200 ;
        RECT  0.685 0.835 0.970 1.180 ;
        RECT  0.650 0.860 0.970 1.180 ;
        RECT  2.080 0.630 2.420 1.180 ;
        RECT  0.650 0.950 2.420 1.180 ;
        RECT  1.575 0.950 1.805 2.490 ;
        RECT  1.575 2.260 2.080 2.490 ;
        RECT  1.850 2.260 2.080 2.830 ;
        RECT  1.850 2.545 2.365 2.830 ;
        RECT  2.680 1.175 3.020 1.515 ;
        RECT  2.680 1.285 3.725 1.515 ;
        RECT  3.495 2.540 4.920 2.900 ;
        RECT  3.495 1.285 3.725 3.100 ;
        RECT  2.760 2.870 3.725 3.100 ;
        RECT  2.760 2.870 3.100 3.880 ;
        RECT  4.900 0.630 5.240 0.950 ;
        RECT  4.900 0.630 5.130 2.310 ;
        RECT  4.900 2.080 5.590 2.310 ;
        RECT  5.180 2.080 5.590 2.455 ;
        RECT  5.180 2.080 5.415 3.360 ;
        RECT  4.230 3.130 5.415 3.360 ;
        RECT  4.230 3.130 4.570 3.840 ;
        RECT  5.360 1.380 6.055 1.720 ;
        RECT  5.820 1.380 6.055 2.480 ;
        RECT  5.820 2.140 7.040 2.480 ;
        RECT  5.820 1.380 6.050 3.880 ;
        RECT  5.670 2.960 6.050 3.880 ;
    END
END NO5I4X2

MACRO NO5I4X1
    CLASS CORE ;
    FOREIGN NO5I4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.955 1.590 4.425 2.110 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 2.860 7.440 3.875 ;
        RECT  7.205 1.360 7.440 3.875 ;
        RECT  6.965 1.360 7.440 1.700 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 1.740 2.690 2.070 ;
        RECT  2.035 1.630 2.405 2.030 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.300 3.265 2.640 ;
        RECT  2.950 2.190 3.265 2.640 ;
        END
    END BN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.320 3.520 1.810 4.020 ;
        END
    END DN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.005 1.290 2.345 ;
        RECT  0.755 2.005 1.135 2.580 ;
        RECT  0.755 2.005 1.110 2.605 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.305 3.505 6.645 5.280 ;
        RECT  4.860 3.615 5.200 5.280 ;
        RECT  3.460 3.910 3.800 5.280 ;
        RECT  2.040 3.060 2.380 5.280 ;
        RECT  1.290 3.060 2.380 3.290 ;
        RECT  1.290 2.750 1.605 3.290 ;
        RECT  1.320 2.720 1.605 3.290 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.225 -0.400 6.565 0.880 ;
        RECT  4.110 -0.400 4.450 0.710 ;
        RECT  1.385 -0.400 1.725 0.710 ;
        RECT  0.180 -0.400 0.520 0.680 ;
        RECT  0.180 -0.400 0.505 0.695 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.410 1.125 1.695 ;
        RECT  0.180 1.410 0.520 4.200 ;
        RECT  0.180 3.860 1.040 4.200 ;
        RECT  0.690 0.835 0.975 1.180 ;
        RECT  0.660 0.865 0.975 1.180 ;
        RECT  2.085 0.630 2.425 1.180 ;
        RECT  0.660 0.950 2.425 1.180 ;
        RECT  1.575 0.950 1.805 2.490 ;
        RECT  1.575 2.260 2.080 2.490 ;
        RECT  1.850 2.260 2.080 2.830 ;
        RECT  1.850 2.545 2.365 2.830 ;
        RECT  2.690 1.185 3.725 1.510 ;
        RECT  3.495 1.185 3.725 3.140 ;
        RECT  3.495 2.640 4.920 2.925 ;
        RECT  2.760 2.910 3.780 3.140 ;
        RECT  2.760 2.910 3.100 3.880 ;
        RECT  4.830 0.745 5.250 1.085 ;
        RECT  4.830 0.745 5.060 2.310 ;
        RECT  4.830 2.015 5.470 2.310 ;
        RECT  5.180 2.015 5.415 3.385 ;
        RECT  4.100 3.155 5.415 3.385 ;
        RECT  4.100 3.155 4.440 3.760 ;
        RECT  5.290 1.445 5.935 1.785 ;
        RECT  5.700 1.445 5.935 2.480 ;
        RECT  5.700 2.140 6.915 2.480 ;
        RECT  5.700 1.445 5.930 3.850 ;
        RECT  5.580 3.550 5.930 3.850 ;
    END
END NO5I4X1

MACRO NO5I4X0
    CLASS CORE ;
    FOREIGN NO5I4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.860 2.395 3.240 ;
        RECT  1.625 2.860 2.395 3.180 ;
        RECT  1.625 2.100 1.965 3.180 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.695 1.030 1.135 1.410 ;
        RECT  0.695 0.630 0.925 1.410 ;
        RECT  0.460 0.630 0.925 0.865 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.583  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.920 3.150 7.385 3.490 ;
        RECT  7.055 1.820 7.385 3.490 ;
        RECT  6.160 1.820 7.385 2.050 ;
        RECT  6.160 0.710 6.390 2.050 ;
        RECT  6.025 0.710 6.390 0.995 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.965 2.250 3.655 2.630 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 1.600 4.235 2.025 ;
        END
    END AN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.295 1.640 3.025 2.020 ;
        RECT  2.295 1.640 2.635 2.310 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.620 -0.400 6.915 1.590 ;
        RECT  4.340 -0.400 4.680 0.790 ;
        RECT  2.180 -0.400 2.520 0.710 ;
        RECT  1.155 -0.400 1.440 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 3.910 6.660 5.280 ;
        RECT  4.920 3.585 5.260 5.280 ;
        RECT  3.420 3.510 3.760 5.280 ;
        RECT  2.070 3.480 2.360 5.280 ;
        RECT  0.980 3.870 1.270 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.095 0.465 3.960 ;
        RECT  0.180 2.045 0.935 2.385 ;
        RECT  0.180 2.045 0.510 3.960 ;
        RECT  1.365 1.020 1.920 1.360 ;
        RECT  1.365 1.020 1.595 1.870 ;
        RECT  0.740 2.830 1.395 3.170 ;
        RECT  1.165 1.640 1.395 3.640 ;
        RECT  1.165 3.410 1.730 3.640 ;
        RECT  1.500 3.410 1.730 4.005 ;
        RECT  1.500 3.665 1.840 4.005 ;
        RECT  3.640 0.655 3.980 1.260 ;
        RECT  3.640 1.030 4.700 1.260 ;
        RECT  4.410 1.030 4.700 1.450 ;
        RECT  4.465 1.030 4.700 2.870 ;
        RECT  3.980 2.530 4.700 2.870 ;
        RECT  3.980 2.530 4.210 3.115 ;
        RECT  2.720 2.885 4.210 3.115 ;
        RECT  2.720 2.885 3.060 3.680 ;
        RECT  4.930 0.710 5.480 0.995 ;
        RECT  4.930 1.975 5.340 2.315 ;
        RECT  4.460 3.125 5.160 3.355 ;
        RECT  4.930 0.710 5.160 3.355 ;
        RECT  4.120 3.345 4.690 3.575 ;
        RECT  4.120 3.345 4.460 3.685 ;
        RECT  5.390 1.405 5.805 1.745 ;
        RECT  5.575 1.405 5.805 3.290 ;
        RECT  5.575 2.600 6.810 2.935 ;
        RECT  5.575 2.600 5.860 3.290 ;
        RECT  5.520 2.950 5.860 3.290 ;
    END
END NO5I4X0

MACRO NO5I3X4
    CLASS CORE ;
    FOREIGN NO5I3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.630 3.450 2.395 3.850 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.138  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.470 3.485 6.950 3.825 ;
        RECT  6.470 2.660 6.700 3.825 ;
        RECT  4.990 1.345 6.650 1.630 ;
        RECT  5.290 2.660 6.700 2.890 ;
        RECT  5.795 1.345 6.175 2.890 ;
        RECT  5.290 2.660 5.630 3.770 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.065 0.525 2.740 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.880 1.315 2.220 ;
        RECT  0.755 1.880 1.135 2.630 ;
        END
    END BN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.295 1.640 8.695 2.220 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.120 8.065 2.630 ;
        RECT  7.390 2.120 8.065 2.460 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.300 2.640 8.640 5.280 ;
        RECT  5.850 4.170 6.190 5.280 ;
        RECT  4.730 4.170 5.070 5.280 ;
        RECT  3.250 3.505 3.590 5.280 ;
        RECT  1.950 4.080 2.290 5.280 ;
        RECT  0.880 3.680 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.125 -0.400 8.470 0.710 ;
        RECT  7.010 -0.400 7.350 0.655 ;
        RECT  5.750 -0.400 6.090 0.655 ;
        RECT  4.230 -0.400 4.570 0.655 ;
        RECT  1.525 -0.400 1.865 0.960 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.095 0.630 2.600 0.940 ;
        RECT  0.225 0.630 0.565 1.440 ;
        RECT  2.095 0.630 2.325 1.440 ;
        RECT  0.225 1.210 2.325 1.440 ;
        RECT  1.390 2.880 1.775 3.220 ;
        RECT  1.545 1.210 1.775 3.220 ;
        RECT  0.290 2.990 1.775 3.220 ;
        RECT  0.290 2.990 0.520 4.215 ;
        RECT  0.180 3.875 0.520 4.215 ;
        RECT  2.555 1.345 3.050 1.685 ;
        RECT  2.710 2.140 3.500 2.480 ;
        RECT  2.710 1.345 3.050 3.170 ;
        RECT  3.040 0.700 3.380 1.040 ;
        RECT  3.040 0.810 3.960 1.040 ;
        RECT  4.830 1.860 5.565 2.200 ;
        RECT  3.730 0.810 3.960 2.940 ;
        RECT  4.830 1.860 5.060 2.940 ;
        RECT  3.730 2.710 5.060 2.940 ;
        RECT  3.970 2.710 4.310 4.180 ;
        RECT  4.300 0.885 7.160 1.115 ;
        RECT  6.930 1.240 7.910 1.580 ;
        RECT  4.300 0.885 4.530 2.480 ;
        RECT  4.190 2.140 4.530 2.480 ;
        RECT  6.930 0.885 7.160 3.135 ;
        RECT  6.930 2.795 7.490 3.135 ;
        RECT  0.225 1.210 1.80 1.440 ;
        RECT  4.300 0.885 6.50 1.115 ;
    END
END NO5I3X4

MACRO NO5I3X2
    CLASS CORE ;
    FOREIGN NO5I3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.420 1.030 3.760 2.035 ;
        RECT  3.275 1.030 3.760 1.410 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.933  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.860 6.870 3.775 ;
        RECT  6.640 1.240 6.870 3.775 ;
        RECT  6.480 1.240 6.870 1.580 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 1.745 2.085 2.070 ;
        RECT  1.385 1.630 1.830 2.020 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.300 2.700 2.640 ;
        RECT  2.320 2.190 2.700 2.640 ;
        END
    END BN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.230 1.245 2.630 ;
        RECT  0.755 2.200 1.215 2.630 ;
        RECT  0.755 2.200 1.000 2.780 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 0.970 1.175 ;
        RECT  0.645 0.850 0.970 1.175 ;
        RECT  0.125 0.885 0.505 1.410 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 4.170 7.380 5.280 ;
        RECT  5.760 2.960 6.100 5.280 ;
        RECT  4.320 3.590 4.660 5.280 ;
        RECT  2.800 3.540 3.140 5.280 ;
        RECT  1.270 2.860 1.570 5.280 ;
        RECT  1.230 2.860 1.570 3.200 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.040 -0.400 7.380 0.720 ;
        RECT  5.920 -0.400 6.260 0.720 ;
        RECT  3.500 -0.400 3.840 0.775 ;
        RECT  1.380 -0.400 1.720 0.955 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.405 1.120 1.870 ;
        RECT  0.180 1.640 1.120 1.870 ;
        RECT  0.180 1.640 0.520 4.230 ;
        RECT  0.180 3.890 1.040 4.230 ;
        RECT  2.080 1.175 2.420 1.515 ;
        RECT  2.080 1.285 3.045 1.515 ;
        RECT  2.815 1.285 3.045 1.935 ;
        RECT  2.930 2.560 4.405 2.900 ;
        RECT  4.080 2.440 4.405 2.900 ;
        RECT  2.930 1.705 3.160 3.100 ;
        RECT  2.135 2.870 3.160 3.100 ;
        RECT  2.135 2.870 2.475 3.210 ;
        RECT  4.270 0.630 4.640 0.950 ;
        RECT  4.270 0.630 4.500 2.210 ;
        RECT  4.270 1.980 5.060 2.210 ;
        RECT  4.635 1.980 5.060 2.455 ;
        RECT  4.635 1.980 4.865 3.360 ;
        RECT  3.600 3.130 4.865 3.360 ;
        RECT  3.600 3.130 3.940 3.840 ;
        RECT  4.730 1.380 5.525 1.720 ;
        RECT  5.290 1.380 5.525 2.480 ;
        RECT  5.290 2.140 6.410 2.480 ;
        RECT  5.095 2.960 5.520 3.880 ;
        RECT  5.290 1.380 5.520 3.880 ;
        RECT  5.040 3.540 5.520 3.880 ;
    END
END NO5I3X2

MACRO NO5I3X1
    CLASS CORE ;
    FOREIGN NO5I3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.400 1.690 3.740 2.030 ;
        RECT  3.400 1.030 3.655 2.030 ;
        RECT  3.275 1.030 3.655 1.410 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 2.860 6.810 3.875 ;
        RECT  6.575 1.230 6.810 3.875 ;
        RECT  6.335 1.230 6.810 1.570 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.910 3.340 2.405 3.850 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.520 2.090 3.025 2.580 ;
        END
    END BN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.150 2.005 1.765 2.580 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.530 0.460 2.240 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.675 3.505 6.015 5.280 ;
        RECT  4.230 3.615 4.570 5.280 ;
        RECT  2.635 3.495 2.975 5.280 ;
        RECT  1.335 2.810 1.680 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.595 -0.400 5.935 1.045 ;
        RECT  3.480 -0.400 3.820 0.710 ;
        RECT  1.585 -0.400 1.925 0.815 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.690 1.070 1.125 1.410 ;
        RECT  0.180 2.815 0.920 3.155 ;
        RECT  0.690 1.070 0.920 4.185 ;
        RECT  0.690 3.845 1.040 4.185 ;
        RECT  2.060 1.170 2.405 1.510 ;
        RECT  2.060 1.170 2.290 3.095 ;
        RECT  3.230 2.690 4.290 2.925 ;
        RECT  3.400 2.640 4.290 2.925 ;
        RECT  2.060 2.810 3.430 3.095 ;
        RECT  4.200 0.745 4.620 1.085 ;
        RECT  4.200 0.745 4.430 2.310 ;
        RECT  4.200 2.015 4.840 2.310 ;
        RECT  4.550 2.015 4.785 3.385 ;
        RECT  3.665 3.155 4.785 3.385 ;
        RECT  3.665 3.155 3.895 3.760 ;
        RECT  3.470 3.420 3.895 3.760 ;
        RECT  4.660 1.445 5.305 1.785 ;
        RECT  5.070 1.445 5.305 2.480 ;
        RECT  5.945 2.140 6.285 2.480 ;
        RECT  5.070 2.250 6.285 2.480 ;
        RECT  5.070 1.445 5.300 3.845 ;
        RECT  4.950 3.550 5.300 3.845 ;
    END
END NO5I3X1

MACRO NO5I3X0
    CLASS CORE ;
    FOREIGN NO5I3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.260 2.860 1.765 3.190 ;
        RECT  1.260 1.800 1.490 3.190 ;
        RECT  0.995 1.800 1.490 2.140 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.155 0.570 3.850 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.584  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 2.250 6.805 2.630 ;
        RECT  6.290 3.170 6.640 3.490 ;
        RECT  6.410 1.820 6.640 3.490 ;
        RECT  5.530 1.820 6.640 2.050 ;
        RECT  5.530 0.710 5.760 2.050 ;
        RECT  5.395 0.710 5.760 0.995 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.335 2.250 3.025 2.580 ;
        RECT  2.335 2.180 2.710 2.580 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.145 1.570 3.605 2.050 ;
        END
    END AN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.720 1.180 2.395 1.410 ;
        RECT  2.015 1.030 2.395 1.410 ;
        RECT  1.720 1.180 2.005 2.310 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.990 -0.400 6.285 1.590 ;
        RECT  3.710 -0.400 4.050 0.790 ;
        RECT  1.550 -0.400 1.890 0.710 ;
        RECT  0.350 -0.400 0.690 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 3.940 6.030 5.280 ;
        RECT  4.365 3.585 4.650 5.280 ;
        RECT  2.790 3.510 3.130 5.280 ;
        RECT  1.440 3.420 1.730 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.535 1.020 1.290 1.360 ;
        RECT  0.535 1.020 0.765 2.925 ;
        RECT  0.185 2.640 0.765 2.925 ;
        RECT  0.185 2.695 1.030 2.925 ;
        RECT  0.800 2.695 1.030 3.905 ;
        RECT  0.800 3.565 1.210 3.905 ;
        RECT  3.010 0.690 3.350 0.975 ;
        RECT  3.120 0.690 3.350 1.340 ;
        RECT  3.120 1.110 4.065 1.340 ;
        RECT  3.255 2.530 4.065 2.870 ;
        RECT  3.835 1.110 4.065 2.870 ;
        RECT  2.090 2.810 3.485 3.040 ;
        RECT  2.090 2.810 2.430 3.680 ;
        RECT  4.300 0.710 4.850 0.995 ;
        RECT  4.300 1.980 4.710 2.265 ;
        RECT  3.905 3.125 4.530 3.355 ;
        RECT  4.300 0.710 4.530 3.355 ;
        RECT  3.490 3.350 4.135 3.650 ;
        RECT  4.760 1.405 5.175 1.745 ;
        RECT  4.945 1.405 5.175 3.290 ;
        RECT  4.945 2.630 6.180 2.965 ;
        RECT  4.890 2.950 5.230 3.290 ;
    END
END NO5I3X0

MACRO NO5I2X4
    CLASS CORE ;
    FOREIGN NO5I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.274  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 1.345 8.695 4.165 ;
        RECT  6.980 2.660 8.695 3.000 ;
        RECT  6.980 1.345 8.695 1.650 ;
        RECT  6.980 2.660 7.320 3.770 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.310 0.525 3.240 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.310 2.650 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.200 2.140 4.915 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.070 3.035 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 1.640 3.755 2.210 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.880 4.210 7.880 5.280 ;
        RECT  6.920 4.170 7.880 5.280 ;
        RECT  6.895 4.190 7.880 5.280 ;
        RECT  4.940 3.780 5.280 5.280 ;
        RECT  2.600 3.615 2.940 5.280 ;
        RECT  1.300 3.650 1.640 5.280 ;
        RECT  0.180 3.650 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.740 -0.400 8.080 0.710 ;
        RECT  6.220 -0.400 6.560 0.770 ;
        RECT  3.680 -0.400 4.020 0.710 ;
        RECT  2.540 -0.400 2.880 0.710 ;
        RECT  1.030 -0.400 1.370 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.640 0.520 0.980 ;
        RECT  0.290 0.640 0.520 2.020 ;
        RECT  0.290 1.790 1.770 2.020 ;
        RECT  1.540 1.880 1.940 2.220 ;
        RECT  1.540 1.790 1.770 3.110 ;
        RECT  0.755 2.880 1.770 3.110 ;
        RECT  0.755 2.880 1.080 3.220 ;
        RECT  1.840 1.235 2.400 1.570 ;
        RECT  1.855 1.235 2.400 1.575 ;
        RECT  5.270 2.140 5.610 2.480 ;
        RECT  2.170 2.860 5.500 3.090 ;
        RECT  5.270 2.140 5.500 3.090 ;
        RECT  2.170 1.235 2.400 3.275 ;
        RECT  2.060 2.935 2.400 3.275 ;
        RECT  3.120 1.110 4.780 1.410 ;
        RECT  4.440 1.110 4.780 1.690 ;
        RECT  4.440 1.460 6.170 1.690 ;
        RECT  5.940 1.880 6.280 2.220 ;
        RECT  5.940 1.460 6.170 3.550 ;
        RECT  4.240 3.320 6.170 3.550 ;
        RECT  4.240 3.320 4.580 4.180 ;
        RECT  5.030 0.700 5.370 1.230 ;
        RECT  5.030 1.000 6.750 1.230 ;
        RECT  6.520 1.880 7.080 2.220 ;
        RECT  6.520 1.000 6.750 4.010 ;
        RECT  5.660 3.780 6.750 4.010 ;
        RECT  5.660 3.780 6.000 4.120 ;
        RECT  2.170 2.860 4.70 3.090 ;
    END
END NO5I2X4

MACRO NO5I2X2
    CLASS CORE ;
    FOREIGN NO5I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.220 2.630 ;
        RECT  0.930 1.750 1.220 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.907  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.850 6.870 3.770 ;
        RECT  6.640 1.240 6.870 3.770 ;
        RECT  6.480 1.240 6.870 1.580 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.305 3.445 1.765 4.015 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.590 0.600 2.050 ;
        RECT  0.115 1.545 0.580 2.050 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.610 3.710 2.595 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.110 2.585 2.630 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 4.170 7.380 5.280 ;
        RECT  5.760 2.960 6.100 5.280 ;
        RECT  4.280 3.840 4.620 5.280 ;
        RECT  3.010 3.935 3.350 5.280 ;
        RECT  1.995 3.595 2.335 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.040 -0.400 7.380 0.720 ;
        RECT  5.920 -0.400 6.260 0.720 ;
        RECT  3.675 -0.400 4.015 0.710 ;
        RECT  1.385 -0.400 1.725 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.085 0.630 2.525 0.955 ;
        RECT  2.085 0.630 2.315 1.430 ;
        RECT  0.785 1.145 2.315 1.430 ;
        RECT  0.800 1.145 1.680 1.475 ;
        RECT  1.450 1.145 1.680 3.100 ;
        RECT  0.795 2.870 1.680 3.100 ;
        RECT  0.180 3.795 0.520 4.140 ;
        RECT  0.180 3.910 1.040 4.140 ;
        RECT  0.795 2.870 1.040 4.250 ;
        RECT  0.685 3.910 1.040 4.250 ;
        RECT  2.685 1.285 3.045 1.625 ;
        RECT  2.450 2.860 3.045 3.195 ;
        RECT  2.815 1.285 3.045 3.705 ;
        RECT  2.815 3.475 4.050 3.705 ;
        RECT  3.710 3.475 4.050 3.900 ;
        RECT  4.475 0.630 4.815 1.145 ;
        RECT  4.270 2.220 4.970 2.560 ;
        RECT  4.270 0.915 4.500 3.245 ;
        RECT  3.715 2.960 4.500 3.245 ;
        RECT  4.730 1.490 5.070 1.830 ;
        RECT  4.730 1.600 5.435 1.830 ;
        RECT  5.200 1.600 5.435 2.540 ;
        RECT  6.070 2.200 6.410 2.540 ;
        RECT  5.200 2.310 6.410 2.540 ;
        RECT  5.200 1.600 5.430 3.880 ;
        RECT  5.040 2.960 5.430 3.880 ;
    END
END NO5I2X2

MACRO NO5I2X1
    CLASS CORE ;
    FOREIGN NO5I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.220 2.630 ;
        RECT  0.930 1.810 1.220 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 2.725 6.810 3.640 ;
        RECT  6.505 1.230 6.810 3.640 ;
        RECT  6.335 1.230 6.810 1.570 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.305 3.445 1.740 4.015 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.605 0.600 2.050 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 1.610 3.780 2.485 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.070 2.635 2.630 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.675 2.780 6.030 5.280 ;
        RECT  3.445 3.845 4.750 5.280 ;
        RECT  1.970 2.860 2.265 5.280 ;
        RECT  1.910 2.860 2.265 3.200 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.595 -0.400 5.935 1.045 ;
        RECT  3.745 -0.400 4.085 0.710 ;
        RECT  1.385 -0.400 1.725 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.085 0.630 2.525 0.955 ;
        RECT  2.085 0.630 2.315 1.430 ;
        RECT  0.800 1.145 2.315 1.430 ;
        RECT  0.800 1.145 1.680 1.485 ;
        RECT  1.450 1.145 1.680 3.100 ;
        RECT  0.795 2.870 1.680 3.100 ;
        RECT  0.180 3.795 1.040 4.140 ;
        RECT  0.795 2.870 1.040 4.250 ;
        RECT  0.685 3.795 1.040 4.250 ;
        RECT  2.755 1.175 3.095 1.515 ;
        RECT  2.865 3.325 4.230 3.615 ;
        RECT  2.865 1.175 3.095 3.865 ;
        RECT  2.640 3.465 3.095 3.865 ;
        RECT  4.545 0.745 4.885 1.150 ;
        RECT  4.195 0.920 4.885 1.150 ;
        RECT  4.195 2.080 4.900 2.420 ;
        RECT  4.195 0.920 4.430 3.065 ;
        RECT  3.650 2.725 4.430 3.065 ;
        RECT  4.660 1.445 5.365 1.785 ;
        RECT  5.130 1.445 5.365 2.480 ;
        RECT  5.130 2.140 6.275 2.480 ;
        RECT  5.130 1.445 5.360 3.130 ;
        RECT  4.970 2.745 5.360 3.130 ;
    END
END NO5I2X1

MACRO NO5I2X0
    CLASS CORE ;
    FOREIGN NO5I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.630 1.205 2.245 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.285 0.570 3.850 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.587  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 3.085 6.805 3.410 ;
        RECT  6.530 1.670 6.805 3.410 ;
        RECT  5.530 1.790 6.805 2.020 ;
        RECT  6.425 1.670 6.805 2.020 ;
        RECT  5.530 0.630 5.760 2.020 ;
        RECT  5.395 0.630 5.760 0.915 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.160 2.250 3.020 2.660 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 1.520 3.605 2.035 ;
        END
    END AN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.805 1.635 2.405 2.020 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.810 3.810 6.150 5.280 ;
        RECT  4.430 3.575 4.770 5.280 ;
        RECT  3.110 3.580 3.450 5.280 ;
        RECT  1.645 3.495 1.985 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.990 -0.400 6.285 1.485 ;
        RECT  5.990 -0.400 6.225 1.550 ;
        RECT  3.795 -0.400 4.130 0.710 ;
        RECT  2.265 -0.400 2.605 0.710 ;
        RECT  0.865 -0.400 1.205 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.565 0.630 1.905 1.170 ;
        RECT  0.180 0.940 1.905 1.170 ;
        RECT  0.180 0.940 0.520 3.045 ;
        RECT  0.180 2.705 1.030 3.045 ;
        RECT  0.800 2.705 1.030 3.985 ;
        RECT  0.800 3.565 1.415 3.985 ;
        RECT  3.095 0.630 3.435 0.915 ;
        RECT  3.205 0.630 3.435 1.260 ;
        RECT  3.205 1.030 4.070 1.260 ;
        RECT  3.780 1.030 4.070 1.370 ;
        RECT  3.835 1.030 4.070 2.495 ;
        RECT  3.250 2.265 4.070 2.495 ;
        RECT  3.250 2.265 3.480 3.280 ;
        RECT  2.345 3.050 3.480 3.280 ;
        RECT  2.345 3.050 2.685 3.845 ;
        RECT  4.595 0.630 4.935 1.095 ;
        RECT  4.300 0.865 4.935 1.095 ;
        RECT  4.300 1.895 4.830 2.235 ;
        RECT  4.300 0.865 4.530 3.200 ;
        RECT  3.710 2.860 4.530 3.200 ;
        RECT  4.760 1.325 5.290 1.665 ;
        RECT  5.060 1.325 5.290 3.210 ;
        RECT  5.060 2.545 6.300 2.880 ;
        RECT  5.010 2.870 5.350 3.210 ;
    END
END NO5I2X0

MACRO NO5I1X4
    CLASS CORE ;
    FOREIGN NO5I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.275 6.820 1.620 ;
        RECT  6.470 2.660 6.810 3.415 ;
        RECT  5.150 2.660 6.810 2.890 ;
        RECT  5.795 1.275 6.175 2.890 ;
        RECT  5.155 1.275 6.820 1.565 ;
        RECT  5.150 2.660 5.490 3.480 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 3.435 0.710 3.855 ;
        END
    END AN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.295 1.030 8.695 2.220 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.140 1.430 2.640 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.407  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.760 1.640 2.395 1.985 ;
        RECT  1.760 1.640 2.375 1.995 ;
        RECT  1.760 1.640 2.100 2.210 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.120 7.605 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.300 2.640 8.640 5.280 ;
        RECT  5.710 4.170 6.050 5.280 ;
        RECT  4.590 4.170 4.930 5.280 ;
        RECT  3.110 3.585 3.450 5.280 ;
        RECT  0.940 3.625 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.295 -0.400 8.640 0.710 ;
        RECT  7.180 -0.400 7.520 0.710 ;
        RECT  5.820 -0.400 6.160 1.045 ;
        RECT  4.450 -0.400 4.790 1.135 ;
        RECT  2.000 -0.400 2.340 0.710 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.175 0.685 0.520 1.040 ;
        RECT  2.490 2.195 2.830 2.680 ;
        RECT  2.525 2.175 2.830 2.680 ;
        RECT  1.840 2.450 2.830 2.680 ;
        RECT  0.290 0.685 0.520 3.100 ;
        RECT  0.180 2.700 0.520 3.100 ;
        RECT  1.840 2.450 2.070 3.100 ;
        RECT  0.180 2.870 2.070 3.100 ;
        RECT  1.440 1.110 2.990 1.410 ;
        RECT  2.760 1.350 3.290 1.690 ;
        RECT  3.060 2.140 3.500 2.480 ;
        RECT  3.060 1.350 3.290 3.250 ;
        RECT  2.570 2.910 3.290 3.250 ;
        RECT  3.300 0.700 3.640 1.040 ;
        RECT  3.300 0.810 3.960 1.040 ;
        RECT  3.730 1.680 4.950 1.910 ;
        RECT  4.750 1.795 5.565 2.025 ;
        RECT  5.225 1.795 5.565 2.225 ;
        RECT  3.730 0.810 3.960 2.940 ;
        RECT  3.830 2.715 4.170 4.180 ;
        RECT  7.740 1.240 8.065 1.580 ;
        RECT  4.210 2.140 4.550 2.485 ;
        RECT  4.540 2.255 4.770 3.940 ;
        RECT  7.150 3.600 8.065 3.830 ;
        RECT  7.835 1.240 8.065 3.830 ;
        RECT  4.540 3.710 7.490 3.940 ;
        RECT  4.540 3.710 6.70 3.940 ;
    END
END NO5I1X4

MACRO NO5I1X2
    CLASS CORE ;
    FOREIGN NO5I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.705 2.050 1.160 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.040 1.115 ;
        RECT  0.750 0.630 1.040 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.770 6.870 3.690 ;
        RECT  6.640 1.240 6.870 3.690 ;
        RECT  6.480 1.240 6.870 1.580 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.765 2.145 4.325 2.630 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.390 2.105 1.775 2.735 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.465 2.860 3.025 3.240 ;
        RECT  2.465 1.975 2.770 3.240 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 4.090 7.380 5.280 ;
        RECT  5.760 2.770 6.100 5.280 ;
        RECT  4.280 3.835 4.620 5.280 ;
        RECT  1.270 3.025 1.555 5.280 ;
        RECT  1.215 3.025 1.555 3.365 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.040 -0.400 7.380 0.720 ;
        RECT  5.920 -0.400 6.260 0.720 ;
        RECT  4.030 -0.400 4.370 0.715 ;
        RECT  2.780 -0.400 3.065 1.470 ;
        RECT  1.380 -0.400 1.720 0.915 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.630 ;
        RECT  0.180 1.590 0.965 1.820 ;
        RECT  0.180 1.590 0.410 4.190 ;
        RECT  0.180 3.850 1.040 4.190 ;
        RECT  0.700 3.850 1.040 4.250 ;
        RECT  4.030 1.175 4.370 1.515 ;
        RECT  3.295 1.285 4.370 1.515 ;
        RECT  3.100 1.815 3.535 2.155 ;
        RECT  3.295 1.285 3.535 3.145 ;
        RECT  3.295 2.860 4.060 3.145 ;
        RECT  2.005 0.630 2.420 0.970 ;
        RECT  4.580 2.090 4.970 2.430 ;
        RECT  2.005 0.630 2.235 3.700 ;
        RECT  3.255 3.375 4.810 3.605 ;
        RECT  4.580 2.090 4.810 3.605 ;
        RECT  2.005 3.470 3.485 3.700 ;
        RECT  2.880 3.470 3.485 3.810 ;
        RECT  4.730 1.170 5.070 1.510 ;
        RECT  4.730 1.280 5.435 1.510 ;
        RECT  5.200 1.280 5.435 2.540 ;
        RECT  6.070 2.200 6.410 2.540 ;
        RECT  5.200 2.310 6.410 2.540 ;
        RECT  5.200 1.280 5.430 3.690 ;
        RECT  5.040 2.770 5.430 3.690 ;
    END
END NO5I1X2

MACRO NO5I1X1
    CLASS CORE ;
    FOREIGN NO5I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.705 2.050 1.160 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.040 1.115 ;
        RECT  0.750 0.630 1.040 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.837  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.250 6.805 2.630 ;
        RECT  6.425 1.075 6.695 2.630 ;
        RECT  6.340 2.760 6.690 3.690 ;
        RECT  6.425 1.075 6.690 3.690 ;
        RECT  6.355 1.075 6.695 1.415 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.765 2.145 4.325 2.580 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.390 2.105 1.775 2.735 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.465 2.860 3.025 3.240 ;
        RECT  2.465 1.975 2.770 3.240 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.745 4.090 6.085 5.280 ;
        RECT  4.265 2.810 4.605 5.280 ;
        RECT  1.270 3.025 1.555 5.280 ;
        RECT  1.215 3.025 1.555 3.365 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.635 -0.400 5.975 1.370 ;
        RECT  3.565 -0.400 3.905 0.655 ;
        RECT  2.780 -0.400 3.065 1.470 ;
        RECT  1.380 -0.400 1.720 0.915 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.630 ;
        RECT  0.180 1.590 0.965 1.820 ;
        RECT  0.180 1.590 0.410 4.190 ;
        RECT  0.180 3.850 1.040 4.190 ;
        RECT  0.700 3.850 1.040 4.250 ;
        RECT  2.005 0.630 2.420 0.970 ;
        RECT  2.005 0.630 2.235 3.820 ;
        RECT  2.005 3.480 3.770 3.820 ;
        RECT  3.430 3.480 3.770 4.010 ;
        RECT  4.360 0.630 4.705 1.115 ;
        RECT  3.295 0.885 4.705 1.115 ;
        RECT  3.180 1.815 3.535 2.155 ;
        RECT  3.295 0.885 3.535 3.150 ;
        RECT  3.295 2.810 3.885 3.150 ;
        RECT  4.405 1.345 5.230 1.655 ;
        RECT  4.985 1.345 5.230 3.110 ;
        RECT  4.985 1.840 6.165 2.180 ;
        RECT  4.985 1.840 5.325 3.110 ;
    END
END NO5I1X1

MACRO NO5I1X0
    CLASS CORE ;
    FOREIGN NO5I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.705 2.050 1.135 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.090 1.115 ;
        RECT  0.750 0.630 1.090 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.345 2.240 6.815 2.640 ;
        RECT  6.345 2.240 6.685 3.050 ;
        RECT  6.345 1.235 6.575 3.050 ;
        RECT  6.040 1.235 6.575 1.560 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.865 1.995 4.325 2.580 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 2.110 1.750 2.745 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.440 2.245 2.980 2.635 ;
        RECT  2.440 1.910 2.725 2.635 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.745 3.505 6.085 5.280 ;
        RECT  4.145 2.810 4.485 5.280 ;
        RECT  1.270 3.575 1.560 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.240 -0.400 5.580 0.985 ;
        RECT  3.410 -0.400 3.755 0.655 ;
        RECT  2.780 -0.400 3.065 1.470 ;
        RECT  1.380 -0.400 1.720 0.905 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.630 ;
        RECT  0.180 1.590 0.965 1.820 ;
        RECT  0.180 1.590 0.410 3.820 ;
        RECT  0.180 3.480 1.040 3.820 ;
        RECT  0.700 3.480 1.040 3.970 ;
        RECT  1.980 0.630 2.420 0.970 ;
        RECT  1.980 0.630 2.210 3.555 ;
        RECT  1.980 3.280 3.505 3.555 ;
        RECT  2.645 3.280 3.505 3.620 ;
        RECT  2.645 3.280 2.985 3.915 ;
        RECT  4.215 0.630 4.555 1.115 ;
        RECT  3.295 0.885 4.555 1.115 ;
        RECT  3.195 1.815 3.535 2.155 ;
        RECT  3.295 0.885 3.535 3.050 ;
        RECT  3.295 2.710 3.670 3.050 ;
        RECT  4.215 1.345 5.230 1.685 ;
        RECT  4.945 1.345 5.230 3.050 ;
        RECT  4.945 1.790 6.105 2.115 ;
        RECT  4.945 1.790 5.285 3.050 ;
    END
END NO5I1X0

MACRO NO4X4
    CLASS CORE ;
    FOREIGN NO4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 1.170 7.385 4.160 ;
        RECT  5.840 2.205 7.385 2.655 ;
        RECT  5.600 3.115 6.070 4.160 ;
        RECT  5.840 1.170 6.070 4.160 ;
        RECT  5.600 1.170 6.070 1.510 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.250 1.135 2.625 ;
        RECT  0.575 1.730 0.890 2.625 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.750 2.250 2.395 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 3.910 3.310 4.250 ;
        RECT  2.645 3.470 3.025 4.250 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.230 1.525 1.765 2.020 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.510 ;
        RECT  4.840 -0.400 5.180 1.000 ;
        RECT  2.990 -0.400 3.330 0.710 ;
        RECT  1.660 -0.400 2.000 0.710 ;
        RECT  0.180 -0.400 0.520 1.040 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 2.920 6.660 5.280 ;
        RECT  4.880 3.180 5.220 5.280 ;
        RECT  3.540 2.720 3.790 5.280 ;
        RECT  3.400 2.720 3.790 3.690 ;
        RECT  1.370 2.865 1.710 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.310 1.400 3.000 1.715 ;
        RECT  2.690 1.400 3.000 3.240 ;
        RECT  2.690 2.150 4.220 2.490 ;
        RECT  2.690 2.150 3.040 3.240 ;
        RECT  0.750 0.940 3.460 1.170 ;
        RECT  0.750 0.940 1.240 1.280 ;
        RECT  0.115 1.270 0.980 1.500 ;
        RECT  3.230 0.940 3.460 1.920 ;
        RECT  3.230 1.690 4.830 1.920 ;
        RECT  4.600 1.690 4.830 2.490 ;
        RECT  4.600 2.150 4.935 2.490 ;
        RECT  0.115 1.270 0.345 4.035 ;
        RECT  0.115 2.865 0.520 4.035 ;
        RECT  3.690 0.700 4.030 1.460 ;
        RECT  3.690 1.230 5.370 1.460 ;
        RECT  5.140 1.230 5.370 2.040 ;
        RECT  5.165 1.890 5.610 2.230 ;
        RECT  5.165 1.890 5.430 2.950 ;
        RECT  4.120 2.720 5.430 2.950 ;
        RECT  4.120 2.720 4.460 4.180 ;
        RECT  0.750 0.940 2.30 1.170 ;
    END
END NO4X4

MACRO NO4X2
    CLASS CORE ;
    FOREIGN NO4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.280  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.045 2.050 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.279  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.315 2.120 1.715 2.685 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.279  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.120 1.085 2.685 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.280  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.160 2.250 5.665 2.770 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.123  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.680 2.250 4.295 2.630 ;
        RECT  3.635 3.025 3.975 3.960 ;
        RECT  3.680 1.680 3.975 3.960 ;
        RECT  3.595 1.680 3.975 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.410 2.985 4.750 5.280 ;
        RECT  2.915 3.080 3.255 5.280 ;
        RECT  1.435 2.990 1.780 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 0.950 ;
        RECT  4.260 -0.400 4.600 0.950 ;
        RECT  1.660 -0.400 2.000 1.350 ;
        RECT  0.180 -0.400 0.520 1.430 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.180 1.240 1.890 ;
        RECT  0.115 1.660 2.270 1.890 ;
        RECT  1.945 1.660 2.270 2.220 ;
        RECT  0.115 1.660 0.345 3.955 ;
        RECT  0.115 2.995 0.625 3.955 ;
        RECT  2.500 0.700 3.220 0.990 ;
        RECT  2.500 0.700 2.730 2.850 ;
        RECT  2.500 2.520 3.450 2.850 ;
        RECT  2.195 2.620 2.535 3.960 ;
        RECT  5.020 1.060 5.360 1.410 ;
        RECT  4.115 1.180 6.125 1.410 ;
        RECT  2.960 1.220 4.305 1.450 ;
        RECT  2.960 1.220 3.300 2.150 ;
        RECT  5.895 1.180 6.125 3.230 ;
        RECT  5.560 3.000 5.900 3.960 ;
        RECT  0.115 1.660 1.20 1.890 ;
        RECT  4.115 1.180 5.60 1.410 ;
    END
END NO4X2

MACRO NO4X1
    CLASS CORE ;
    FOREIGN NO4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.760 1.640 5.100 1.980 ;
        RECT  3.905 1.640 5.100 1.875 ;
        RECT  3.905 1.030 4.285 1.875 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.950 1.775 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.150 1.135 3.240 ;
        RECT  0.700 2.150 1.135 2.490 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.186  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.250 5.725 2.630 ;
        RECT  5.440 1.670 5.725 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.210 1.030 3.025 1.420 ;
        RECT  2.450 2.645 2.790 3.565 ;
        RECT  2.210 2.645 2.790 2.875 ;
        RECT  2.210 1.030 2.440 2.875 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.690 3.670 5.030 5.280 ;
        RECT  3.170 2.645 3.510 5.280 ;
        RECT  1.610 2.870 1.955 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.470 -0.400 6.010 0.710 ;
        RECT  0.350 -0.400 1.965 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.185 1.170 1.365 1.510 ;
        RECT  0.185 1.170 0.465 3.940 ;
        RECT  0.185 2.815 0.525 3.940 ;
        RECT  0.185 3.600 0.610 3.940 ;
        RECT  3.295 1.070 3.620 2.335 ;
        RECT  2.690 1.995 3.620 2.335 ;
        RECT  2.690 2.105 4.270 2.335 ;
        RECT  3.930 2.105 4.270 3.065 ;
        RECT  5.070 1.070 6.185 1.410 ;
        RECT  5.955 1.070 6.185 3.200 ;
        RECT  5.680 2.860 6.185 3.200 ;
        RECT  5.680 2.860 5.910 4.250 ;
        RECT  5.320 3.910 5.910 4.250 ;
    END
END NO4X1

MACRO NO4X0
    CLASS CORE ;
    FOREIGN NO4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.760 1.615 5.100 1.930 ;
        RECT  3.905 1.615 5.100 1.875 ;
        RECT  3.905 1.030 4.285 1.875 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.250 5.725 2.630 ;
        RECT  5.440 1.670 5.725 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.055 1.765 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.480 1.135 3.240 ;
        RECT  0.700 2.480 1.135 2.820 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.170 1.030 3.025 1.510 ;
        RECT  2.350 2.615 2.690 3.200 ;
        RECT  2.170 1.030 2.400 2.845 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.750 3.510 5.090 5.280 ;
        RECT  3.150 2.860 3.490 5.280 ;
        RECT  1.650 3.040 1.995 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.470 -0.400 6.010 0.710 ;
        RECT  0.425 -0.400 1.965 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 1.365 1.510 ;
        RECT  0.180 1.170 0.465 3.940 ;
        RECT  0.180 3.040 0.520 3.940 ;
        RECT  0.180 3.600 0.610 3.940 ;
        RECT  3.255 1.070 3.580 2.335 ;
        RECT  2.630 1.995 3.580 2.335 ;
        RECT  2.630 2.105 4.290 2.335 ;
        RECT  3.950 2.105 4.290 3.200 ;
        RECT  5.070 1.070 6.185 1.385 ;
        RECT  5.955 1.070 6.185 3.200 ;
        RECT  5.780 2.860 6.010 4.130 ;
        RECT  5.320 3.790 6.010 4.130 ;
    END
END NO4X0

MACRO NO4I3X4
    CLASS CORE ;
    FOREIGN NO4I3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.355 0.570 3.920 ;
        END
    END CN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.765 3.430 2.125 ;
        RECT  2.645 1.635 3.030 2.125 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.955 2.810 4.480 3.275 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.230 2.095 1.765 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.002  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.760 2.860 9.270 3.265 ;
        RECT  8.900 1.270 9.270 3.265 ;
        RECT  7.720 1.270 9.270 1.610 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.320 3.565 8.660 5.280 ;
        RECT  7.050 3.560 7.425 5.280 ;
        RECT  5.570 2.780 5.910 5.280 ;
        RECT  4.260 3.815 4.600 5.280 ;
        RECT  2.780 3.510 3.120 5.280 ;
        RECT  0.940 2.885 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.295 -0.400 8.635 1.035 ;
        RECT  7.025 -0.400 7.365 1.040 ;
        RECT  4.445 -0.400 4.785 1.515 ;
        RECT  2.545 -0.400 2.885 1.180 ;
        RECT  0.940 -0.400 1.285 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.975 0.630 2.315 1.170 ;
        RECT  0.180 0.940 2.315 1.170 ;
        RECT  0.180 0.705 0.520 2.980 ;
        RECT  1.740 1.400 2.340 1.695 ;
        RECT  2.110 1.400 2.340 2.980 ;
        RECT  2.110 2.580 3.010 2.920 ;
        RECT  2.110 2.580 2.480 2.980 ;
        RECT  3.290 1.175 4.105 1.515 ;
        RECT  3.875 1.745 5.000 2.085 ;
        RECT  3.875 1.175 4.105 2.580 ;
        RECT  3.495 2.350 4.105 2.580 ;
        RECT  3.495 2.350 3.725 3.880 ;
        RECT  3.495 3.535 3.840 3.880 ;
        RECT  5.155 1.070 5.510 1.410 ;
        RECT  5.235 1.070 5.510 2.450 ;
        RECT  5.235 2.110 7.070 2.450 ;
        RECT  4.795 2.315 5.465 2.545 ;
        RECT  4.795 2.315 5.135 3.560 ;
        RECT  5.875 0.700 6.215 1.880 ;
        RECT  5.875 1.650 7.490 1.880 ;
        RECT  7.300 1.855 8.670 2.195 ;
        RECT  7.300 1.745 7.530 2.910 ;
        RECT  6.335 2.680 7.530 2.910 ;
        RECT  6.335 2.680 6.675 4.160 ;
        RECT  0.180 0.940 1.80 1.170 ;
    END
END NO4I3X4

MACRO NO4I3X2
    CLASS CORE ;
    FOREIGN NO4I3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.320 3.520 1.810 4.020 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.930 2.860 7.435 3.240 ;
        RECT  7.150 1.245 7.380 3.240 ;
        RECT  6.930 2.745 7.285 3.665 ;
        RECT  6.910 1.245 7.380 1.585 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 1.740 2.635 2.125 ;
        RECT  2.015 1.635 2.400 2.025 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 2.130 3.820 2.640 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.940 1.290 2.280 ;
        RECT  0.755 1.940 1.135 2.580 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.665 2.745 7.990 5.280 ;
        RECT  6.400 4.115 6.740 5.280 ;
        RECT  4.885 2.745 5.225 5.280 ;
        RECT  3.520 3.810 3.860 5.280 ;
        RECT  2.040 3.060 2.380 5.280 ;
        RECT  1.320 3.060 2.380 3.290 ;
        RECT  1.320 2.720 1.605 3.290 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.650 -0.400 7.995 1.585 ;
        RECT  6.380 -0.400 6.720 0.710 ;
        RECT  3.680 -0.400 4.020 0.775 ;
        RECT  1.385 -0.400 1.725 0.710 ;
        RECT  0.180 -0.400 0.520 0.680 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.410 1.125 1.695 ;
        RECT  0.180 1.410 0.520 4.150 ;
        RECT  0.180 3.810 1.040 4.150 ;
        RECT  0.635 0.890 0.975 1.180 ;
        RECT  2.085 0.630 2.425 1.180 ;
        RECT  0.635 0.950 2.425 1.180 ;
        RECT  1.555 0.950 1.785 2.490 ;
        RECT  1.555 2.260 2.080 2.490 ;
        RECT  1.850 2.260 2.080 2.830 ;
        RECT  1.850 2.545 2.365 2.830 ;
        RECT  2.690 1.175 3.095 1.515 ;
        RECT  2.865 1.175 3.095 3.825 ;
        RECT  2.865 3.350 4.655 3.580 ;
        RECT  4.325 3.350 4.655 3.690 ;
        RECT  2.760 3.460 3.100 3.825 ;
        RECT  4.470 1.155 4.825 2.365 ;
        RECT  4.470 2.025 5.720 2.365 ;
        RECT  4.245 2.035 4.475 3.110 ;
        RECT  4.085 2.770 4.475 3.110 ;
        RECT  5.180 1.225 5.520 1.585 ;
        RECT  5.180 1.355 6.245 1.585 ;
        RECT  6.010 1.355 6.245 2.480 ;
        RECT  6.010 2.140 6.920 2.480 ;
        RECT  6.010 1.355 6.240 2.975 ;
        RECT  5.605 2.745 6.240 2.975 ;
        RECT  5.605 2.745 5.945 3.665 ;
    END
END NO4I3X2

MACRO NO4I3X1
    CLASS CORE ;
    FOREIGN NO4I3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.320 3.520 1.810 4.020 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 2.745 6.805 3.665 ;
        RECT  6.575 1.245 6.805 3.665 ;
        RECT  6.335 1.245 6.805 1.585 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 1.740 2.635 2.125 ;
        RECT  2.015 1.635 2.400 2.025 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 1.925 3.635 2.635 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.940 1.290 2.280 ;
        RECT  0.755 1.940 1.135 2.580 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.880 4.065 6.220 5.280 ;
        RECT  4.575 3.590 4.915 5.280 ;
        RECT  3.520 3.910 3.860 5.280 ;
        RECT  2.040 3.060 2.380 5.280 ;
        RECT  1.320 3.060 2.380 3.290 ;
        RECT  1.320 2.720 1.605 3.290 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.595 -0.400 5.935 1.045 ;
        RECT  3.680 -0.400 4.020 0.710 ;
        RECT  1.385 -0.400 1.725 0.710 ;
        RECT  0.180 -0.400 0.520 0.690 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.410 1.125 1.695 ;
        RECT  0.180 1.410 0.520 4.150 ;
        RECT  0.180 3.810 1.040 4.150 ;
        RECT  0.635 0.890 0.975 1.180 ;
        RECT  2.085 0.630 2.425 1.180 ;
        RECT  0.635 0.950 2.425 1.180 ;
        RECT  1.555 0.950 1.785 2.490 ;
        RECT  1.555 2.260 2.080 2.490 ;
        RECT  1.850 2.260 2.080 2.830 ;
        RECT  1.850 2.545 2.365 2.830 ;
        RECT  2.690 1.175 3.095 1.515 ;
        RECT  2.865 1.175 3.095 3.850 ;
        RECT  2.865 3.350 4.345 3.660 ;
        RECT  4.015 3.350 4.345 3.690 ;
        RECT  2.760 3.510 3.100 3.850 ;
        RECT  4.470 0.745 4.825 1.090 ;
        RECT  4.200 0.860 4.825 1.090 ;
        RECT  4.200 2.025 5.145 2.365 ;
        RECT  4.200 0.860 4.430 3.110 ;
        RECT  3.765 2.825 4.430 3.110 ;
        RECT  4.660 1.445 4.945 1.785 ;
        RECT  4.660 1.555 5.670 1.785 ;
        RECT  5.435 1.555 5.670 2.480 ;
        RECT  5.435 2.140 6.345 2.480 ;
        RECT  5.435 1.555 5.665 3.120 ;
        RECT  5.085 2.760 5.665 3.120 ;
    END
END NO4I3X1

MACRO NO4I3X0
    CLASS CORE ;
    FOREIGN NO4I3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.040 2.260 2.380 2.740 ;
        RECT  2.040 1.960 2.345 2.740 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.695 1.030 1.135 1.410 ;
        RECT  0.695 0.630 0.925 1.410 ;
        RECT  0.460 0.630 0.925 0.915 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.558  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.110 2.765 6.805 3.240 ;
        RECT  6.575 0.630 6.805 3.240 ;
        RECT  6.410 0.630 6.805 0.970 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.210 2.150 3.605 2.670 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.590 1.470 3.020 2.020 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.510 3.560 5.850 5.280 ;
        RECT  3.910 3.390 4.270 5.280 ;
        RECT  2.180 3.410 2.520 5.280 ;
        RECT  0.980 3.370 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.660 -0.400 6.000 0.715 ;
        RECT  4.140 -0.400 4.480 0.710 ;
        RECT  2.510 -0.400 2.850 0.915 ;
        RECT  1.155 -0.400 1.495 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.160 0.465 3.620 ;
        RECT  0.180 2.100 1.350 2.425 ;
        RECT  0.180 2.100 0.520 3.620 ;
        RECT  1.580 1.160 1.920 1.500 ;
        RECT  1.070 2.685 1.810 3.010 ;
        RECT  1.580 1.160 1.810 3.900 ;
        RECT  1.580 3.560 1.950 3.900 ;
        RECT  3.340 0.630 3.910 0.915 ;
        RECT  3.680 0.630 3.910 1.920 ;
        RECT  3.835 1.690 4.205 2.030 ;
        RECT  3.835 1.690 4.065 3.130 ;
        RECT  2.880 2.900 4.065 3.130 ;
        RECT  2.880 2.900 3.220 3.710 ;
        RECT  4.140 1.170 4.665 1.455 ;
        RECT  4.435 1.805 4.925 2.145 ;
        RECT  4.435 1.170 4.665 2.860 ;
        RECT  4.295 2.520 4.665 2.860 ;
        RECT  4.840 0.630 5.385 0.970 ;
        RECT  5.155 2.220 6.290 2.535 ;
        RECT  5.155 0.630 5.385 3.350 ;
        RECT  4.710 3.090 5.385 3.350 ;
        RECT  4.710 3.090 5.050 3.710 ;
    END
END NO4I3X0

MACRO NO4I2X4
    CLASS CORE ;
    FOREIGN NO4I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.002  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.130 2.860 8.640 3.265 ;
        RECT  8.275 1.265 8.640 3.265 ;
        RECT  8.270 1.305 8.640 3.265 ;
        RECT  7.090 1.305 8.640 1.610 ;
        RECT  7.090 1.265 7.375 1.610 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.765 2.800 2.125 ;
        RECT  2.015 1.635 2.400 2.125 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 2.810 3.850 3.275 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.600 2.120 1.135 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 0.940 1.685 1.170 ;
        RECT  1.345 0.630 1.685 1.170 ;
        RECT  0.115 0.940 0.570 1.420 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.665 -0.400 8.005 1.045 ;
        RECT  6.395 -0.400 6.735 1.040 ;
        RECT  3.815 -0.400 4.155 1.515 ;
        RECT  1.915 -0.400 2.255 1.405 ;
        RECT  0.310 -0.400 0.655 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.690 3.565 8.030 5.280 ;
        RECT  6.420 3.560 6.795 5.280 ;
        RECT  4.940 2.795 5.280 5.280 ;
        RECT  3.630 3.815 3.970 5.280 ;
        RECT  2.150 3.510 2.490 5.280 ;
        RECT  0.310 2.885 0.650 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.110 1.400 1.685 1.695 ;
        RECT  1.455 1.400 1.685 2.980 ;
        RECT  1.455 2.580 2.380 2.980 ;
        RECT  2.660 1.175 3.260 1.515 ;
        RECT  3.030 1.790 4.370 2.130 ;
        RECT  3.030 1.175 3.260 2.580 ;
        RECT  2.865 2.350 3.095 3.880 ;
        RECT  2.865 3.535 3.210 3.880 ;
        RECT  4.525 1.055 4.880 1.395 ;
        RECT  4.605 1.055 4.880 2.450 ;
        RECT  4.605 2.110 6.440 2.450 ;
        RECT  4.165 2.360 4.835 2.590 ;
        RECT  4.165 2.360 4.505 3.560 ;
        RECT  5.245 0.700 5.585 1.880 ;
        RECT  5.245 1.650 6.860 1.880 ;
        RECT  6.670 1.750 6.905 2.230 ;
        RECT  6.670 1.890 8.040 2.230 ;
        RECT  6.670 1.750 6.900 2.925 ;
        RECT  5.705 2.680 6.900 2.925 ;
        RECT  5.705 2.680 6.045 4.160 ;
    END
END NO4I2X4

MACRO NO4I2X2
    CLASS CORE ;
    FOREIGN NO4I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.300 2.860 6.790 3.240 ;
        RECT  6.520 1.240 6.750 3.240 ;
        RECT  6.300 2.745 6.640 3.665 ;
        RECT  6.280 1.240 6.750 1.580 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.700 1.740 2.005 2.465 ;
        RECT  1.385 1.635 1.770 1.970 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.695 2.110 3.135 2.665 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.175 1.275 2.660 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.950 0.990 1.180 ;
        RECT  0.635 0.875 0.990 1.180 ;
        RECT  0.125 0.950 0.550 1.375 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.020 -0.400 7.365 1.580 ;
        RECT  5.750 -0.400 6.090 0.710 ;
        RECT  3.080 -0.400 3.420 0.710 ;
        RECT  1.385 -0.400 1.725 0.955 ;
        RECT  0.180 -0.400 0.520 0.675 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.020 2.745 7.360 5.280 ;
        RECT  5.770 4.065 6.110 5.280 ;
        RECT  4.255 2.745 4.595 5.280 ;
        RECT  2.890 3.810 3.230 5.280 ;
        RECT  1.370 2.890 1.710 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.785 1.410 1.125 1.890 ;
        RECT  0.180 1.605 1.125 1.890 ;
        RECT  0.180 1.605 0.520 4.150 ;
        RECT  0.180 3.810 1.040 4.150 ;
        RECT  2.090 1.175 2.465 1.515 ;
        RECT  2.235 1.175 2.465 3.845 ;
        RECT  2.235 3.350 4.025 3.580 ;
        RECT  3.695 3.350 4.025 3.690 ;
        RECT  2.130 3.505 2.470 3.845 ;
        RECT  3.770 0.710 4.125 2.365 ;
        RECT  3.770 2.025 5.090 2.365 ;
        RECT  3.455 2.035 3.795 3.110 ;
        RECT  4.550 1.200 4.890 1.560 ;
        RECT  4.550 1.330 5.615 1.560 ;
        RECT  5.380 1.330 5.615 2.480 ;
        RECT  5.380 2.140 6.290 2.480 ;
        RECT  5.380 1.330 5.610 2.975 ;
        RECT  4.975 2.745 5.610 2.975 ;
        RECT  4.975 2.745 5.315 3.665 ;
    END
END NO4I2X2

MACRO NO4I2X1
    CLASS CORE ;
    FOREIGN NO4I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.745 6.175 3.665 ;
        RECT  5.945 1.250 6.175 3.665 ;
        RECT  5.705 1.250 6.175 1.590 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.720 1.690 2.005 2.460 ;
        RECT  1.385 1.640 1.765 2.020 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.695 1.925 3.010 2.630 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.230 1.290 2.630 ;
        RECT  0.750 2.210 1.255 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.950 0.975 1.180 ;
        RECT  0.635 0.875 0.975 1.180 ;
        RECT  0.125 0.950 0.505 1.370 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.220 4.065 5.560 5.280 ;
        RECT  3.950 3.590 4.290 5.280 ;
        RECT  2.890 3.910 3.230 5.280 ;
        RECT  1.410 2.860 1.750 5.280 ;
        RECT  1.240 2.860 1.750 3.210 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.965 -0.400 5.305 1.045 ;
        RECT  3.080 -0.400 3.420 0.710 ;
        RECT  1.385 -0.400 1.725 0.800 ;
        RECT  0.180 -0.400 0.520 0.675 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.765 1.410 1.125 1.830 ;
        RECT  0.180 1.600 1.125 1.830 ;
        RECT  0.180 1.600 0.520 4.205 ;
        RECT  0.180 3.865 1.040 4.205 ;
        RECT  2.090 1.175 2.465 1.460 ;
        RECT  2.235 1.175 2.465 3.830 ;
        RECT  2.235 3.350 3.720 3.635 ;
        RECT  3.375 3.350 3.720 3.690 ;
        RECT  2.130 3.490 2.470 3.830 ;
        RECT  3.870 0.745 4.225 1.125 ;
        RECT  3.570 0.895 4.225 1.125 ;
        RECT  3.570 2.025 4.515 2.365 ;
        RECT  3.570 0.895 3.800 3.110 ;
        RECT  3.135 2.825 3.800 3.110 ;
        RECT  4.030 1.445 4.315 1.785 ;
        RECT  4.030 1.555 5.040 1.785 ;
        RECT  4.805 1.555 5.040 2.480 ;
        RECT  4.805 2.140 5.715 2.480 ;
        RECT  4.805 1.555 5.035 3.120 ;
        RECT  4.455 2.780 5.035 3.120 ;
    END
END NO4I2X1

MACRO NO4I2X0
    CLASS CORE ;
    FOREIGN NO4I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.410 2.250 1.850 2.715 ;
        RECT  1.410 2.210 1.805 2.715 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.540 0.720 2.030 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.558  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.480 2.765 6.175 3.240 ;
        RECT  5.945 0.630 6.175 3.240 ;
        RECT  5.780 0.630 6.175 0.970 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 2.260 2.975 2.630 ;
        RECT  2.620 2.140 2.975 2.630 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.960 1.485 2.390 2.035 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.880 3.560 5.220 5.280 ;
        RECT  3.280 3.360 3.620 5.280 ;
        RECT  1.555 3.400 1.895 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.030 -0.400 5.370 0.975 ;
        RECT  3.510 -0.400 3.850 0.710 ;
        RECT  1.880 -0.400 2.220 0.960 ;
        RECT  0.350 -0.400 0.690 0.865 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.950 1.160 1.290 1.500 ;
        RECT  0.405 2.640 1.180 2.980 ;
        RECT  0.950 1.160 1.180 3.890 ;
        RECT  0.950 3.550 1.320 3.890 ;
        RECT  2.710 0.630 3.280 0.960 ;
        RECT  3.050 0.630 3.280 1.920 ;
        RECT  3.205 1.690 3.575 2.030 ;
        RECT  3.205 1.690 3.435 3.130 ;
        RECT  2.250 2.900 3.435 3.130 ;
        RECT  2.250 2.900 2.590 3.700 ;
        RECT  3.510 1.170 4.035 1.455 ;
        RECT  3.805 1.805 4.295 2.145 ;
        RECT  3.805 1.170 4.035 2.880 ;
        RECT  3.665 2.540 4.035 2.880 ;
        RECT  4.210 0.630 4.755 0.970 ;
        RECT  4.525 2.220 5.660 2.535 ;
        RECT  4.525 0.630 4.755 3.365 ;
        RECT  4.080 3.135 4.755 3.365 ;
        RECT  4.080 3.135 4.420 3.680 ;
    END
END NO4I2X0

MACRO NO4I1X4
    CLASS CORE ;
    FOREIGN NO4I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.356  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.845 1.785 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.356  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.525 0.505 2.295 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 2.845 8.695 3.900 ;
        RECT  8.300 1.110 8.640 3.900 ;
        RECT  7.035 2.030 8.640 2.260 ;
        RECT  7.035 1.075 7.265 2.860 ;
        RECT  6.860 2.660 7.205 3.900 ;
        RECT  6.860 1.075 7.265 1.415 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 3.450 4.350 3.980 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.356  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.445 2.400 2.045 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.575 2.660 7.920 5.280 ;
        RECT  6.100 3.080 6.440 5.280 ;
        RECT  4.580 2.640 4.920 5.280 ;
        RECT  1.850 2.860 2.190 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.450 ;
        RECT  6.100 -0.400 6.440 1.285 ;
        RECT  3.370 -0.400 3.710 0.670 ;
        RECT  1.885 -0.400 2.225 1.145 ;
        RECT  0.445 -0.400 0.785 1.155 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.165 0.875 1.505 1.615 ;
        RECT  0.735 1.385 1.505 1.615 ;
        RECT  0.735 1.385 0.965 2.870 ;
        RECT  0.515 2.640 0.855 4.250 ;
        RECT  0.165 3.965 0.855 4.250 ;
        RECT  3.970 1.360 4.275 2.375 ;
        RECT  3.090 2.120 4.160 2.460 ;
        RECT  3.820 2.120 4.160 3.005 ;
        RECT  2.605 0.805 2.945 1.130 ;
        RECT  2.605 0.900 4.735 1.130 ;
        RECT  4.505 0.900 4.735 2.390 ;
        RECT  4.505 2.050 6.160 2.390 ;
        RECT  2.630 0.805 2.860 3.135 ;
        RECT  2.630 2.795 3.340 3.135 ;
        RECT  3.000 2.795 3.340 3.885 ;
        RECT  4.965 0.700 5.250 1.745 ;
        RECT  4.965 1.515 6.630 1.745 ;
        RECT  6.400 2.045 6.805 2.385 ;
        RECT  6.400 1.515 6.630 2.850 ;
        RECT  5.340 2.620 6.630 2.850 ;
        RECT  5.340 2.620 5.680 4.160 ;
        RECT  2.605 0.900 3.90 1.130 ;
    END
END NO4I1X4

MACRO NO4I1X2
    CLASS CORE ;
    FOREIGN NO4I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.050 1.155 3.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.040 1.115 ;
        RECT  0.750 0.630 1.040 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.495 1.225 6.805 3.250 ;
        RECT  6.320 2.660 6.665 3.550 ;
        RECT  6.320 1.225 6.805 1.565 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.900 3.400 2.240 ;
        RECT  2.645 1.640 3.035 2.240 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.075 1.810 2.710 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.035 2.660 7.380 5.280 ;
        RECT  5.600 2.640 5.940 5.280 ;
        RECT  4.160 2.640 4.500 5.280 ;
        RECT  1.420 3.290 1.760 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.040 -0.400 7.380 1.585 ;
        RECT  5.560 -0.400 5.900 1.695 ;
        RECT  2.780 -0.400 3.120 0.690 ;
        RECT  1.380 -0.400 1.720 0.890 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.820 ;
        RECT  0.180 1.590 1.120 1.820 ;
        RECT  0.180 1.590 0.410 4.175 ;
        RECT  0.180 3.835 0.520 4.175 ;
        RECT  0.180 3.890 1.040 4.175 ;
        RECT  0.700 3.890 1.040 4.250 ;
        RECT  3.380 1.380 3.860 1.670 ;
        RECT  3.630 1.380 3.860 2.995 ;
        RECT  2.500 2.655 3.860 2.995 ;
        RECT  2.040 0.630 2.420 1.150 ;
        RECT  3.660 0.805 4.000 1.150 ;
        RECT  2.040 0.920 4.000 1.150 ;
        RECT  2.040 0.630 2.270 3.665 ;
        RECT  2.040 3.325 2.910 3.665 ;
        RECT  4.330 0.880 4.670 2.275 ;
        RECT  4.330 2.045 6.265 2.275 ;
        RECT  4.880 2.045 6.265 2.385 ;
        RECT  4.880 2.045 5.220 3.560 ;
    END
END NO4I1X2

MACRO NO4I1X1
    CLASS CORE ;
    FOREIGN NO4I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.050 1.155 3.240 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.040 1.115 ;
        RECT  0.750 0.630 1.040 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.955 1.225 6.185 3.250 ;
        RECT  5.675 2.660 6.020 3.550 ;
        RECT  5.780 1.225 6.185 1.565 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.980 1.845 3.400 2.130 ;
        RECT  2.645 1.640 3.145 2.020 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.075 1.770 2.710 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.115 3.940 5.455 5.280 ;
        RECT  3.635 2.890 3.975 5.280 ;
        RECT  1.270 3.455 1.560 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.020 -0.400 5.360 0.875 ;
        RECT  2.780 -0.400 3.120 0.690 ;
        RECT  1.380 -0.400 1.720 0.885 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.820 ;
        RECT  0.180 1.590 1.120 1.820 ;
        RECT  0.180 1.590 0.410 4.175 ;
        RECT  0.180 3.835 1.040 4.175 ;
        RECT  0.700 3.835 1.040 4.250 ;
        RECT  3.380 1.380 3.860 1.615 ;
        RECT  3.630 1.380 3.860 2.590 ;
        RECT  2.460 2.360 3.860 2.590 ;
        RECT  2.460 2.360 3.255 2.700 ;
        RECT  2.915 2.360 3.255 3.190 ;
        RECT  2.000 0.630 2.420 1.150 ;
        RECT  3.660 0.805 4.000 1.150 ;
        RECT  2.000 0.920 4.000 1.150 ;
        RECT  2.000 0.630 2.230 3.955 ;
        RECT  2.000 3.615 2.750 3.955 ;
        RECT  4.230 0.630 4.530 2.275 ;
        RECT  4.355 2.045 5.725 2.385 ;
        RECT  4.355 2.045 4.695 3.200 ;
        RECT  2.000 0.920 3.50 1.150 ;
    END
END NO4I1X1

MACRO NO4I1X0
    CLASS CORE ;
    FOREIGN NO4I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.050 1.135 3.250 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.885 1.040 1.115 ;
        RECT  0.750 0.630 1.040 1.115 ;
        RECT  0.125 0.885 0.505 1.360 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.558  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.715 2.710 6.185 3.245 ;
        RECT  5.955 0.630 6.185 3.245 ;
        RECT  5.780 0.630 6.185 0.970 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.955 1.895 3.390 2.235 ;
        RECT  2.645 1.640 3.150 2.020 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 2.075 1.750 2.710 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.115 3.455 5.455 5.280 ;
        RECT  2.915 3.315 3.855 5.280 ;
        RECT  1.270 3.480 1.610 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.040 -0.400 5.380 0.965 ;
        RECT  2.780 -0.400 3.120 0.690 ;
        RECT  1.380 -0.400 1.720 0.920 ;
        RECT  0.180 -0.400 0.520 0.655 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 1.345 1.120 1.820 ;
        RECT  0.180 1.590 1.120 1.820 ;
        RECT  0.180 1.590 0.410 3.865 ;
        RECT  0.180 3.525 1.040 3.865 ;
        RECT  0.700 3.525 1.040 3.960 ;
        RECT  3.380 1.380 3.905 1.665 ;
        RECT  2.440 2.300 2.725 2.695 ;
        RECT  2.440 2.465 3.905 2.695 ;
        RECT  3.620 1.380 3.905 2.945 ;
        RECT  3.515 2.465 3.905 2.945 ;
        RECT  1.980 0.630 2.420 1.150 ;
        RECT  3.660 0.805 4.000 1.150 ;
        RECT  1.980 0.920 4.000 1.150 ;
        RECT  1.980 0.630 2.210 3.810 ;
        RECT  1.980 3.470 2.555 3.810 ;
        RECT  4.230 0.630 4.600 0.990 ;
        RECT  4.315 0.630 4.600 3.520 ;
        RECT  4.315 2.065 5.725 2.405 ;
        RECT  4.315 2.065 4.655 3.520 ;
        RECT  1.980 0.920 3.60 1.150 ;
    END
END NO4I1X0

MACRO NO3X4
    CLASS CORE ;
    FOREIGN NO3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.642  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.945 2.250 6.935 2.480 ;
        RECT  6.595 2.120 6.935 2.480 ;
        RECT  4.775 2.120 5.115 2.480 ;
        RECT  2.945 2.120 3.290 2.480 ;
        RECT  1.200 2.860 3.175 3.090 ;
        RECT  2.945 2.120 3.175 3.090 ;
        RECT  1.200 2.860 1.765 3.240 ;
        RECT  1.200 2.120 1.430 3.240 ;
        RECT  1.090 2.120 1.430 2.460 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.642  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.765 2.120 2.585 2.630 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.649  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.265 1.640 7.615 2.210 ;
        RECT  0.125 1.640 7.615 1.890 ;
        RECT  3.620 1.640 4.445 2.020 ;
        RECT  0.125 1.640 0.760 2.210 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.031  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.405 2.710 8.075 2.940 ;
        RECT  7.845 1.180 8.075 2.940 ;
        RECT  0.900 1.180 8.075 1.410 ;
        RECT  6.990 1.050 7.330 1.410 ;
        RECT  5.685 2.710 6.025 4.180 ;
        RECT  5.460 1.050 5.800 1.410 ;
        RECT  3.905 1.030 4.285 1.410 ;
        RECT  2.000 3.320 3.635 3.550 ;
        RECT  3.405 2.710 3.635 3.550 ;
        RECT  2.420 1.050 2.760 1.410 ;
        RECT  2.000 3.320 2.340 4.180 ;
        RECT  0.900 1.050 1.240 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.620 3.240 7.960 5.280 ;
        RECT  3.865 3.170 4.205 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 0.710 ;
        RECT  6.230 -0.400 6.570 0.950 ;
        RECT  4.700 -0.400 5.040 0.950 ;
        RECT  3.180 -0.400 3.520 0.950 ;
        RECT  1.660 -0.400 2.000 0.950 ;
        RECT  0.180 -0.400 0.520 1.390 ;
        END
    END gnd!
END NO3X4

MACRO NO3X2
    CLASS CORE ;
    FOREIGN NO3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.440 2.120 3.785 2.460 ;
        RECT  1.735 2.860 3.670 3.090 ;
        RECT  3.440 2.120 3.670 3.090 ;
        RECT  1.735 2.120 1.965 3.090 ;
        RECT  1.385 2.120 1.965 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.575 2.120 3.115 2.630 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.115 1.640 4.455 2.220 ;
        RECT  0.705 1.640 4.455 1.890 ;
        RECT  0.705 1.640 1.135 2.210 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.043  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.680 4.915 2.910 ;
        RECT  4.685 1.030 4.915 2.910 ;
        RECT  0.900 1.180 4.915 1.410 ;
        RECT  3.905 1.030 4.915 1.410 ;
        RECT  2.535 3.320 4.130 3.550 ;
        RECT  3.900 2.680 4.130 3.550 ;
        RECT  2.535 3.320 2.875 4.180 ;
        RECT  2.420 1.050 2.760 1.410 ;
        RECT  0.900 1.050 1.240 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.360 3.140 4.700 5.280 ;
        RECT  0.715 2.690 1.055 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.520 -0.400 4.860 0.710 ;
        RECT  3.290 -0.400 3.635 0.710 ;
        RECT  1.660 -0.400 2.000 0.950 ;
        RECT  0.180 -0.400 0.520 1.390 ;
        END
    END gnd!
END NO3X2

MACRO NO3X1
    CLASS CORE ;
    FOREIGN NO3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.690 1.480 2.030 ;
        RECT  0.755 1.690 1.145 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.830 1.510 2.415 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.525 2.460 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.451  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 0.940 3.035 1.410 ;
        RECT  2.060 2.640 2.875 2.980 ;
        RECT  2.645 0.940 2.875 2.980 ;
        RECT  2.420 0.700 2.760 1.280 ;
        RECT  0.900 0.940 3.035 1.280 ;
        RECT  2.060 2.640 2.400 4.180 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.430 2.900 0.770 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.660 -0.400 2.000 0.710 ;
        RECT  0.180 -0.400 0.520 1.115 ;
        END
    END gnd!
END NO3X1

MACRO NO3X0
    CLASS CORE ;
    FOREIGN NO3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.071  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.810 3.480 2.405 3.860 ;
        RECT  2.175 0.630 2.405 3.860 ;
        RECT  0.700 1.170 2.405 1.510 ;
        RECT  2.000 0.630 2.405 1.510 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.510 2.210 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.160 1.320 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.855 1.930 3.250 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.180 3.465 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.530 -0.400 1.640 0.710 ;
        END
    END gnd!
END NO3X0

MACRO NO3I2X4
    CLASS CORE ;
    FOREIGN NO3I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.640  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.065 1.375 8.405 2.220 ;
        RECT  7.275 1.375 8.405 1.605 ;
        RECT  5.350 1.215 7.495 1.445 ;
        RECT  1.195 1.655 5.580 1.895 ;
        RECT  5.350 1.215 5.580 1.895 ;
        RECT  4.420 1.655 5.245 2.020 ;
        RECT  1.195 1.655 1.535 2.220 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.362  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.475 3.155 9.965 3.385 ;
        RECT  9.735 0.900 9.965 3.385 ;
        RECT  7.715 0.900 9.965 1.130 ;
        RECT  8.475 2.910 8.705 3.385 ;
        RECT  5.810 2.910 8.705 3.140 ;
        RECT  7.715 0.755 8.055 1.145 ;
        RECT  4.780 0.755 8.055 0.985 ;
        RECT  6.485 2.910 6.825 4.180 ;
        RECT  6.230 0.645 6.570 0.985 ;
        RECT  2.800 2.710 6.040 2.940 ;
        RECT  1.675 1.185 5.120 1.425 ;
        RECT  4.780 0.755 5.120 1.425 ;
        RECT  3.220 1.030 3.655 1.425 ;
        RECT  2.800 2.710 3.140 4.180 ;
        RECT  1.675 1.050 2.015 1.425 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.465 3.620 9.805 3.960 ;
        RECT  7.685 3.620 9.805 3.850 ;
        RECT  7.685 3.470 8.065 3.850 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.060 0.505 2.630 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.345 4.080 8.685 5.280 ;
        RECT  4.665 3.170 5.005 5.280 ;
        RECT  0.930 3.320 1.270 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.460 -0.400 8.800 0.670 ;
        RECT  3.980 -0.400 4.320 0.955 ;
        RECT  2.445 -0.400 2.785 0.955 ;
        RECT  0.955 -0.400 1.295 1.370 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.700 0.520 1.830 ;
        RECT  0.180 1.600 0.965 1.830 ;
        RECT  5.810 1.675 7.055 1.905 ;
        RECT  6.835 1.835 7.735 2.085 ;
        RECT  7.395 1.835 7.735 2.170 ;
        RECT  1.865 2.125 2.205 2.480 ;
        RECT  3.745 2.125 4.090 2.480 ;
        RECT  5.575 2.125 6.040 2.480 ;
        RECT  1.865 2.250 6.040 2.480 ;
        RECT  5.810 1.675 6.040 2.480 ;
        RECT  0.735 2.450 2.095 2.680 ;
        RECT  0.735 1.600 0.965 3.090 ;
        RECT  0.180 2.860 0.965 3.090 ;
        RECT  0.180 2.860 0.520 4.180 ;
        RECT  6.270 2.135 6.610 2.680 ;
        RECT  6.270 2.450 9.505 2.680 ;
        RECT  9.220 1.360 9.505 2.925 ;
        RECT  9.105 2.450 9.505 2.925 ;
        RECT  1.865 2.250 5.70 2.480 ;
        RECT  6.270 2.450 8.60 2.680 ;
    END
END NO3I2X4

MACRO NO3I2X2
    CLASS CORE ;
    FOREIGN NO3I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.095 0.570 2.630 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.020 1.640 6.345 2.220 ;
        RECT  2.680 1.640 6.345 1.890 ;
        RECT  4.535 1.640 4.915 2.000 ;
        RECT  2.680 1.640 3.020 2.400 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.957  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.440 2.690 6.805 2.920 ;
        RECT  6.575 1.030 6.805 2.920 ;
        RECT  2.920 1.180 6.805 1.410 ;
        RECT  5.795 1.030 6.805 1.410 ;
        RECT  4.440 2.690 4.780 4.180 ;
        RECT  4.440 1.120 4.780 1.410 ;
        RECT  2.920 1.120 3.260 1.410 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.260 2.120 1.765 2.630 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.265 3.150 6.605 5.280 ;
        RECT  2.605 3.090 2.945 5.280 ;
        RECT  0.940 3.320 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 0.710 ;
        RECT  5.195 -0.400 5.540 0.710 ;
        RECT  3.680 -0.400 4.020 0.950 ;
        RECT  2.200 1.120 2.540 1.430 ;
        RECT  2.260 -0.400 2.540 1.430 ;
        RECT  0.940 -0.400 1.280 0.670 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.690 0.630 2.030 0.940 ;
        RECT  0.800 0.900 1.920 1.130 ;
        RECT  0.180 1.240 1.030 1.580 ;
        RECT  0.800 0.900 1.030 3.090 ;
        RECT  0.180 2.860 1.030 3.090 ;
        RECT  0.180 2.860 0.520 3.200 ;
        RECT  1.500 1.360 1.840 1.890 ;
        RECT  1.500 1.660 2.225 1.890 ;
        RECT  3.515 2.120 3.855 2.460 ;
        RECT  5.345 2.120 5.690 2.460 ;
        RECT  3.515 2.230 5.690 2.460 ;
        RECT  3.515 2.120 3.745 2.860 ;
        RECT  1.995 2.630 3.745 2.860 ;
        RECT  1.995 1.660 2.225 3.250 ;
        RECT  1.685 2.910 2.225 3.250 ;
        RECT  3.515 2.230 4.90 2.460 ;
    END
END NO3I2X2

MACRO NO3I2X1
    CLASS CORE ;
    FOREIGN NO3I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.780 1.515 2.160 ;
        RECT  0.755 1.640 1.510 2.160 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.456  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 1.220 3.215 1.560 ;
        RECT  2.630 2.630 3.025 4.180 ;
        RECT  2.630 1.015 2.860 4.180 ;
        RECT  1.540 1.015 2.860 1.245 ;
        RECT  1.540 0.905 1.880 1.245 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.390 0.820 3.850 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.035 4.295 2.640 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.330 3.670 3.670 5.280 ;
        RECT  1.050 2.850 1.390 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.625 -0.400 3.965 0.900 ;
        RECT  2.300 -0.400 2.640 0.710 ;
        RECT  0.780 -0.400 1.120 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.300 0.525 1.640 ;
        RECT  0.220 1.300 0.525 2.980 ;
        RECT  1.845 1.645 2.185 2.620 ;
        RECT  0.220 2.390 2.185 2.620 ;
        RECT  0.220 2.390 0.560 2.980 ;
        RECT  3.445 1.360 3.965 1.705 ;
        RECT  3.090 1.935 3.675 2.275 ;
        RECT  3.445 1.360 3.675 3.210 ;
        RECT  3.445 2.870 4.230 3.210 ;
    END
END NO3I2X1

MACRO NO3I2X0
    CLASS CORE ;
    FOREIGN NO3I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.971  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.020 2.710 3.330 3.045 ;
        RECT  2.020 2.250 2.395 3.045 ;
        RECT  2.020 0.630 2.250 3.045 ;
        RECT  1.725 0.630 2.250 0.970 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.390 1.625 1.790 2.200 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.040 1.145 2.620 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.700 1.615 4.285 2.020 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  2.990 3.560 3.330 5.280 ;
        RECT  1.410 2.635 1.750 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.250 -0.400 3.590 0.710 ;
        RECT  2.480 -0.400 2.790 1.640 ;
        RECT  1.025 -0.400 1.365 1.005 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.290 1.300 0.765 1.640 ;
        RECT  0.290 2.850 0.950 3.140 ;
        RECT  0.290 1.300 0.525 3.145 ;
        RECT  0.460 2.850 0.800 3.700 ;
        RECT  3.850 0.910 4.190 1.250 ;
        RECT  3.240 0.965 4.190 1.250 ;
        RECT  3.240 0.965 3.470 2.480 ;
        RECT  2.750 1.920 3.470 2.260 ;
        RECT  3.235 2.250 4.130 2.480 ;
        RECT  3.790 2.250 4.130 3.700 ;
    END
END NO3I2X0

MACRO NO3I1X4
    CLASS CORE ;
    FOREIGN NO3I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.640  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.435 1.880 7.775 2.220 ;
        RECT  7.435 1.375 7.665 2.220 ;
        RECT  6.645 1.375 7.665 1.605 ;
        RECT  4.720 1.215 6.865 1.445 ;
        RECT  0.515 1.655 4.950 1.895 ;
        RECT  4.720 1.215 4.950 1.895 ;
        RECT  3.790 1.655 4.615 2.020 ;
        RECT  0.515 1.655 0.855 2.220 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.362  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.015 3.155 9.335 3.385 ;
        RECT  9.105 0.900 9.335 3.385 ;
        RECT  7.085 0.900 9.335 1.130 ;
        RECT  8.015 2.910 8.245 3.385 ;
        RECT  5.180 2.910 8.245 3.140 ;
        RECT  7.085 0.755 7.425 1.145 ;
        RECT  4.150 0.755 7.425 0.985 ;
        RECT  5.855 2.910 6.195 4.180 ;
        RECT  5.600 0.645 5.940 0.985 ;
        RECT  2.170 2.710 5.410 2.940 ;
        RECT  0.995 1.185 4.490 1.425 ;
        RECT  4.150 0.755 4.490 1.425 ;
        RECT  2.590 1.030 3.025 1.425 ;
        RECT  2.170 2.710 2.510 4.180 ;
        RECT  0.995 1.050 1.335 1.425 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.486  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.835 3.620 9.175 3.960 ;
        RECT  7.055 3.620 9.175 3.850 ;
        RECT  7.055 3.470 7.435 3.850 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.642  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.765 1.835 7.105 2.170 ;
        RECT  6.205 1.835 7.105 2.065 ;
        RECT  5.180 1.675 6.425 1.905 ;
        RECT  1.235 2.250 5.410 2.480 ;
        RECT  5.180 1.675 5.410 2.480 ;
        RECT  4.945 2.125 5.410 2.480 ;
        RECT  3.115 2.125 3.460 2.480 ;
        RECT  1.235 2.250 1.765 2.630 ;
        RECT  1.235 2.125 1.575 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.715 4.080 8.055 5.280 ;
        RECT  4.035 3.170 4.375 5.280 ;
        RECT  0.275 2.640 0.615 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.830 -0.400 8.170 0.670 ;
        RECT  3.350 -0.400 3.690 0.955 ;
        RECT  1.815 -0.400 2.155 0.955 ;
        RECT  0.235 -0.400 0.575 1.425 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  5.640 2.135 5.980 2.680 ;
        RECT  5.640 2.450 8.875 2.680 ;
        RECT  8.590 1.360 8.875 2.925 ;
        RECT  8.475 2.450 8.875 2.925 ;
        RECT  5.640 2.450 7.70 2.680 ;
    END
END NO3I1X4

MACRO NO3I1X2
    CLASS CORE ;
    FOREIGN NO3I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.120 0.620 2.630 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.730 1.640 5.070 2.220 ;
        RECT  1.310 1.640 5.070 1.890 ;
        RECT  1.310 1.640 1.765 2.020 ;
        RECT  1.310 1.640 1.650 2.400 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.944  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.020 2.860 5.545 3.090 ;
        RECT  5.315 1.030 5.545 3.090 ;
        RECT  1.500 1.180 5.545 1.410 ;
        RECT  4.540 1.030 5.545 1.410 ;
        RECT  3.020 2.860 3.360 4.180 ;
        RECT  3.020 1.120 3.360 1.410 ;
        RECT  1.500 1.120 1.840 1.410 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.821  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.120 4.400 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.970 3.320 5.310 5.280 ;
        RECT  1.070 3.325 1.410 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.100 -0.400 5.440 0.710 ;
        RECT  3.780 -0.400 4.120 0.950 ;
        RECT  2.260 -0.400 2.600 0.950 ;
        RECT  0.740 -0.400 1.080 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.240 1.080 1.580 ;
        RECT  2.560 2.120 3.600 2.460 ;
        RECT  0.850 1.240 1.080 3.095 ;
        RECT  0.310 2.860 1.080 3.095 ;
        RECT  2.560 2.120 2.790 3.095 ;
        RECT  0.310 2.865 2.790 3.095 ;
        RECT  0.310 2.860 0.650 3.200 ;
        RECT  0.310 2.865 1.60 3.095 ;
    END
END NO3I1X2

MACRO NO3I1X1
    CLASS CORE ;
    FOREIGN NO3I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.835 1.560 2.395 1.970 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.412  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.110 1.560 2.450 ;
        RECT  0.755 2.110 1.145 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.456  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.660 3.425 2.890 ;
        RECT  3.160 1.100 3.425 2.890 ;
        RECT  3.085 1.100 3.425 1.560 ;
        RECT  1.700 1.100 3.425 1.330 ;
        RECT  2.630 2.660 3.025 4.180 ;
        RECT  1.700 0.990 2.040 1.330 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.450 0.805 3.855 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.050 3.355 1.390 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.460 -0.400 2.800 0.710 ;
        RECT  0.980 -0.400 1.320 1.315 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.065 0.520 1.410 ;
        RECT  2.615 2.110 2.930 2.430 ;
        RECT  1.920 2.200 2.930 2.430 ;
        RECT  0.280 1.065 0.520 3.205 ;
        RECT  1.920 2.200 2.150 3.090 ;
        RECT  0.280 2.860 2.150 3.090 ;
        RECT  0.280 2.860 0.620 3.205 ;
    END
END NO3I1X1

MACRO NO3I1X0
    CLASS CORE ;
    FOREIGN NO3I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.996  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 3.065 2.940 3.405 ;
        RECT  2.015 3.065 2.395 3.850 ;
        RECT  1.655 3.065 2.940 3.350 ;
        RECT  1.655 0.710 1.885 3.350 ;
        RECT  1.480 0.710 1.885 1.050 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.860 1.425 3.190 ;
        RECT  1.195 2.480 1.425 3.190 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.450 0.505 2.170 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.900 3.025 2.630 ;
        RECT  2.115 1.900 3.025 2.240 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.980 3.420 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.180 -0.400 2.520 1.550 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.935 0.520 1.220 ;
        RECT  0.180 0.990 0.965 1.220 ;
        RECT  0.735 0.990 0.965 2.630 ;
        RECT  0.180 2.400 0.965 2.630 ;
        RECT  0.180 2.400 0.520 4.120 ;
    END
END NO3I1X0

MACRO NO2X4
    CLASS CORE ;
    FOREIGN NO2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.938  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.180 1.400 4.430 3.110 ;
        RECT  3.850 2.900 4.295 4.180 ;
        RECT  3.975 1.400 4.430 1.690 ;
        RECT  1.480 2.900 4.295 3.130 ;
        RECT  0.940 1.400 2.800 1.690 ;
        RECT  1.810 1.400 2.040 3.130 ;
        RECT  1.480 2.860 1.820 4.180 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.750 0.940 5.100 2.630 ;
        RECT  0.290 0.940 5.100 1.170 ;
        RECT  2.940 1.875 3.305 2.210 ;
        RECT  3.045 0.940 3.305 2.210 ;
        RECT  0.125 1.640 0.520 2.220 ;
        RECT  0.290 0.940 0.520 2.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.601  LAYER MET1  ;
        ANTENNAGATEAREA 1.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.270 2.440 3.950 2.670 ;
        RECT  3.610 2.330 3.950 2.670 ;
        RECT  2.270 1.920 2.610 2.670 ;
        RECT  0.755 2.250 1.580 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.000 2.860 5.340 5.280 ;
        RECT  2.700 3.370 3.040 5.280 ;
        RECT  0.330 2.860 0.670 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  0.180 -0.400 5.080 0.710 ;
        END
    END gnd!
END NO2X4

MACRO NO2X2
    CLASS CORE ;
    FOREIGN NO2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.469  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.400 2.410 1.690 ;
        RECT  1.385 2.860 1.780 4.180 ;
        RECT  1.550 1.400 1.780 4.180 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.742  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.300 2.075 2.870 2.415 ;
        RECT  2.640 0.940 2.870 2.415 ;
        RECT  0.280 0.940 2.870 1.170 ;
        RECT  0.125 1.625 0.510 2.220 ;
        RECT  0.280 0.940 0.510 2.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.742  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.320 2.630 ;
        RECT  0.980 1.920 1.320 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.550 2.860 2.890 5.280 ;
        RECT  0.250 2.860 0.590 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  0.180 -0.400 2.970 0.710 ;
        END
    END gnd!
END NO2X2

MACRO NO2X1
    CLASS CORE ;
    FOREIGN NO2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.061  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.330 2.860 1.775 4.180 ;
        RECT  1.545 1.210 1.775 4.180 ;
        RECT  0.780 1.210 1.775 1.550 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.625 0.520 2.265 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.315 2.630 ;
        RECT  1.030 1.940 1.315 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  0.180 2.850 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  0.180 -0.400 1.710 0.710 ;
        END
    END gnd!
END NO2X1

MACRO NO2X0
    CLASS CORE ;
    FOREIGN NO2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.611  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.330 2.860 1.775 3.310 ;
        RECT  1.545 1.170 1.775 3.310 ;
        RECT  0.950 1.170 1.775 1.510 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.475 0.595 2.030 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.315 2.630 ;
        RECT  0.975 2.020 1.315 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  0.180 2.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  0.180 -0.400 1.290 0.710 ;
        END
    END gnd!
END NO2X0

MACRO NO2I1X4
    CLASS CORE ;
    FOREIGN NO2I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.630  LAYER MET1  ;
        ANTENNAGATEAREA 1.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.150 2.440 4.960 2.670 ;
        RECT  4.620 2.330 4.960 2.670 ;
        RECT  3.150 1.920 3.490 2.670 ;
        RECT  1.995 2.055 2.405 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.938  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.900 5.440 3.130 ;
        RECT  5.190 1.400 5.440 3.130 ;
        RECT  4.905 1.400 5.440 1.690 ;
        RECT  4.535 2.900 4.970 4.180 ;
        RECT  1.870 1.400 3.730 1.690 ;
        RECT  2.330 2.860 2.920 3.130 ;
        RECT  2.690 1.400 2.920 3.130 ;
        RECT  2.330 2.860 2.670 4.180 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.484  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.685 0.940 2.220 ;
        END
    END AN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  1.110 -0.400 6.010 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 2.910 6.120 5.280 ;
        RECT  3.480 3.370 3.820 5.280 ;
        RECT  1.180 2.910 1.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.350 0.940 6.020 1.170 ;
        RECT  0.350 0.700 0.700 1.455 ;
        RECT  3.960 0.940 4.210 2.210 ;
        RECT  3.870 1.875 4.210 2.210 ;
        RECT  1.410 1.970 1.760 2.310 ;
        RECT  1.410 0.940 1.640 2.680 ;
        RECT  0.460 2.450 1.640 2.680 ;
        RECT  5.670 0.940 6.020 2.680 ;
        RECT  0.460 2.450 0.800 4.180 ;
        RECT  0.350 0.940 5.70 1.170 ;
    END
END NO2I1X4

MACRO NO2I1X2
    CLASS CORE ;
    FOREIGN NO2I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.742  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.685 2.630 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.705 2.095 1.155 2.630 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.469  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.865 1.400 3.535 1.690 ;
        RECT  2.475 2.860 3.145 3.250 ;
        RECT  2.915 1.400 3.145 3.250 ;
        RECT  2.475 2.860 2.815 4.180 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.625 2.860 3.965 5.280 ;
        RECT  1.325 2.860 1.665 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.305 -0.400 4.095 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.405 0.940 3.995 1.170 ;
        RECT  0.235 1.200 1.635 1.545 ;
        RECT  1.405 0.940 1.635 2.270 ;
        RECT  1.385 1.200 1.635 2.270 ;
        RECT  1.385 1.920 1.725 2.270 ;
        RECT  3.765 0.940 3.995 2.385 ;
        RECT  3.665 2.045 3.995 2.385 ;
        RECT  0.235 1.200 0.475 3.200 ;
        RECT  0.235 2.860 0.925 3.200 ;
        RECT  0.565 2.860 0.925 3.780 ;
        RECT  1.405 0.940 2.60 1.170 ;
    END
END NO2I1X2

MACRO NO2I1X1
    CLASS CORE ;
    FOREIGN NO2I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.028  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.175 1.030 2.405 3.005 ;
        RECT  2.000 2.720 2.340 4.010 ;
        RECT  1.430 1.240 2.405 1.580 ;
        RECT  2.015 1.030 2.405 1.580 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.371  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 1.880 1.300 2.215 ;
        RECT  0.750 1.610 1.135 2.215 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.415 0.605 3.910 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.850 3.670 1.190 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  2.000 -0.400 2.340 0.710 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.965 ;
        RECT  1.540 1.890 1.945 2.230 ;
        RECT  1.540 1.890 1.770 2.675 ;
        RECT  0.290 2.445 1.770 2.675 ;
        RECT  0.290 0.630 0.520 3.185 ;
        RECT  0.180 2.845 0.520 3.185 ;
    END
END NO2I1X1

MACRO NO2I1X0
    CLASS CORE ;
    FOREIGN NO2I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.616  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 1.165 2.395 3.225 ;
        RECT  2.015 1.030 2.395 3.225 ;
        RECT  1.470 1.165 2.395 1.505 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.164  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.195 2.250 1.765 2.630 ;
        RECT  1.195 1.890 1.540 2.630 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.555 0.505 2.120 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.810 3.535 1.150 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.170 ;
        RECT  0.180 0.940 0.965 1.170 ;
        RECT  0.735 0.940 0.965 3.215 ;
        RECT  0.180 2.890 0.965 3.215 ;
        RECT  0.180 2.985 1.695 3.215 ;
        RECT  1.465 2.985 1.695 3.885 ;
        RECT  1.465 3.540 2.100 3.885 ;
    END
END NO2I1X0

MACRO NA8X1
    CLASS CORE ;
    FOREIGN NA8X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.070 0.535 2.655 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.455 3.820 8.065 4.160 ;
        RECT  7.685 3.470 8.065 4.160 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.735 2.100 6.175 2.670 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.405 2.330 6.805 3.190 ;
        END
    END E
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 2.000 2.630 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END G
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.995 1.995 8.695 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.865 3.470 9.325 4.215 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.859  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.275 1.500 5.560 1.840 ;
        RECT  4.745 2.860 5.545 3.190 ;
        RECT  4.745 2.850 5.505 3.190 ;
        RECT  5.275 1.500 5.505 3.190 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.295 3.825 8.635 5.280 ;
        RECT  6.745 3.880 7.090 5.280 ;
        RECT  5.345 4.170 5.685 5.280 ;
        RECT  2.180 4.020 2.520 5.280 ;
        RECT  0.780 3.680 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  6.935 -0.400 7.275 1.410 ;
        RECT  3.240 1.430 4.585 1.770 ;
        RECT  3.240 -0.400 3.580 1.770 ;
        RECT  1.640 -0.400 1.980 0.960 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  2.230 1.260 2.500 3.145 ;
        RECT  0.180 2.885 2.500 3.145 ;
        RECT  0.180 2.885 1.710 3.200 ;
        RECT  1.480 2.885 1.710 4.020 ;
        RECT  1.480 3.680 1.820 4.020 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  4.040 0.630 5.045 0.970 ;
        RECT  2.780 0.630 3.010 2.375 ;
        RECT  2.780 2.090 5.045 2.375 ;
        RECT  4.815 0.630 5.045 2.430 ;
        RECT  3.600 2.090 5.045 2.430 ;
        RECT  3.600 2.090 3.940 3.195 ;
        RECT  5.705 0.800 6.270 1.140 ;
        RECT  6.040 0.800 6.270 1.870 ;
        RECT  6.040 1.640 7.265 1.870 ;
        RECT  7.035 1.640 7.265 3.650 ;
        RECT  3.990 3.420 7.265 3.650 ;
        RECT  3.990 3.420 4.330 3.795 ;
        RECT  6.045 3.420 6.385 4.010 ;
        RECT  8.595 1.130 9.085 1.470 ;
        RECT  8.745 0.630 9.085 1.470 ;
        RECT  9.040 1.185 9.270 3.235 ;
        RECT  7.505 2.895 9.270 3.235 ;
        RECT  0.290 1.590 1.80 1.820 ;
        RECT  0.180 2.885 1.30 3.145 ;
        RECT  2.780 2.090 4.40 2.375 ;
        RECT  3.990 3.420 6.60 3.650 ;
    END
END NA8X1

MACRO NA8X0
    CLASS CORE ;
    FOREIGN NA8X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.530 2.655 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.215 2.095 8.065 2.435 ;
        RECT  7.685 1.640 8.065 2.435 ;
        END
    END B
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 1.360 ;
        END
    END G
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 1.990 2.335 ;
        RECT  1.385 2.050 1.765 2.630 ;
        END
    END H
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.830 2.330 6.175 3.195 ;
        RECT  5.795 2.330 6.175 3.190 ;
        RECT  5.775 2.330 6.175 2.670 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.105 2.100 5.545 2.670 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.785 0.810 7.435 1.410 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.421  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.645 1.500 4.930 1.840 ;
        RECT  4.535 2.860 4.915 3.275 ;
        RECT  4.140 2.850 4.875 3.190 ;
        RECT  4.645 1.500 4.875 3.275 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.225 3.280 8.695 3.850 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.195 -0.400 6.535 1.410 ;
        RECT  3.240 1.430 3.955 1.770 ;
        RECT  3.240 -0.400 3.580 1.770 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.410 3.500 7.750 5.280 ;
        RECT  6.140 3.965 6.480 5.280 ;
        RECT  4.740 3.965 5.080 5.280 ;
        RECT  2.180 3.510 2.520 5.280 ;
        RECT  0.780 3.510 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  2.220 1.260 2.500 3.145 ;
        RECT  0.180 2.885 2.500 3.145 ;
        RECT  0.180 2.885 1.820 3.200 ;
        RECT  1.480 2.885 1.820 3.740 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  4.040 0.630 4.415 0.970 ;
        RECT  2.780 0.630 3.010 2.235 ;
        RECT  4.080 1.965 4.415 2.290 ;
        RECT  2.780 2.005 4.415 2.235 ;
        RECT  4.185 0.630 4.415 2.290 ;
        RECT  3.425 2.005 4.415 2.290 ;
        RECT  3.425 2.005 3.655 3.850 ;
        RECT  3.425 3.510 3.765 3.850 ;
        RECT  4.810 0.800 5.640 1.140 ;
        RECT  5.410 0.800 5.640 1.870 ;
        RECT  5.410 1.640 6.635 1.870 ;
        RECT  5.440 3.420 5.780 3.735 ;
        RECT  6.405 1.640 6.635 3.735 ;
        RECT  3.995 3.505 6.635 3.735 ;
        RECT  3.995 3.505 4.330 3.850 ;
        RECT  8.265 0.630 8.655 1.470 ;
        RECT  8.210 2.650 8.655 2.990 ;
        RECT  8.315 0.630 8.655 2.990 ;
        RECT  6.865 2.705 8.655 2.990 ;
        RECT  6.865 2.705 7.150 3.190 ;
        RECT  0.290 1.590 1.70 1.820 ;
        RECT  0.180 2.885 1.60 3.145 ;
        RECT  3.995 3.505 5.60 3.735 ;
    END
END NA8X0

MACRO NA7X1
    CLASS CORE ;
    FOREIGN NA7X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.070 0.535 2.655 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.310 3.220 8.700 3.855 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.735 2.100 6.175 2.670 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.405 2.330 6.805 3.190 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.495 2.095 8.065 2.435 ;
        RECT  7.685 1.690 8.065 2.435 ;
        RECT  7.685 1.665 8.040 2.435 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.859  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.275 1.500 5.560 1.840 ;
        RECT  4.745 2.860 5.545 3.190 ;
        RECT  4.745 2.850 5.505 3.190 ;
        RECT  5.275 1.500 5.505 3.190 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 2.000 2.630 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.935 -0.400 7.275 1.410 ;
        RECT  3.240 1.430 4.585 1.770 ;
        RECT  3.240 -0.400 3.580 1.770 ;
        RECT  1.640 -0.400 1.980 0.960 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.745 3.880 7.990 5.280 ;
        RECT  7.650 3.825 7.990 5.280 ;
        RECT  5.345 4.170 5.685 5.280 ;
        RECT  2.180 4.020 2.520 5.280 ;
        RECT  0.780 3.685 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.315 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  2.230 1.315 2.500 3.145 ;
        RECT  0.180 2.885 2.500 3.145 ;
        RECT  0.180 2.885 1.710 3.200 ;
        RECT  1.480 2.885 1.710 4.020 ;
        RECT  1.480 3.680 1.820 4.020 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  4.040 0.630 5.045 0.970 ;
        RECT  2.780 0.630 3.010 2.375 ;
        RECT  2.780 2.090 5.045 2.375 ;
        RECT  4.815 0.630 5.045 2.430 ;
        RECT  3.600 2.090 5.045 2.430 ;
        RECT  3.600 2.090 3.940 3.195 ;
        RECT  5.705 0.800 6.270 1.140 ;
        RECT  6.040 0.800 6.270 1.870 ;
        RECT  6.040 1.640 7.265 1.870 ;
        RECT  7.035 1.640 7.265 3.650 ;
        RECT  3.990 3.420 7.265 3.650 ;
        RECT  3.990 3.420 4.330 3.850 ;
        RECT  6.045 3.420 6.385 4.010 ;
        RECT  8.165 0.630 8.655 0.915 ;
        RECT  8.165 0.630 8.550 1.470 ;
        RECT  8.320 0.630 8.550 2.990 ;
        RECT  7.495 2.760 8.550 2.990 ;
        RECT  7.495 2.760 7.800 3.190 ;
        RECT  0.290 1.590 1.90 1.820 ;
        RECT  0.180 2.885 1.70 3.145 ;
        RECT  2.780 2.090 4.00 2.375 ;
        RECT  3.990 3.420 6.30 3.650 ;
    END
END NA7X1

MACRO NA7X0
    CLASS CORE ;
    FOREIGN NA7X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.530 2.655 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 3.220 8.065 3.850 ;
        RECT  7.540 3.220 8.065 3.565 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 1.360 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 2.000 2.630 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.330 6.175 3.190 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.105 2.100 5.545 2.670 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.865 2.095 7.435 2.435 ;
        RECT  7.055 1.690 7.435 2.435 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.421  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.645 1.500 4.930 1.840 ;
        RECT  4.140 2.860 4.915 3.190 ;
        RECT  4.140 2.850 4.875 3.190 ;
        RECT  4.645 1.500 4.875 3.190 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.040 -0.400 6.380 1.410 ;
        RECT  3.240 1.430 3.955 1.770 ;
        RECT  3.240 -0.400 3.580 1.770 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.140 3.880 7.360 5.280 ;
        RECT  7.020 3.825 7.360 5.280 ;
        RECT  4.740 3.880 5.080 5.280 ;
        RECT  2.180 3.510 2.520 5.280 ;
        RECT  0.780 3.510 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  2.230 1.260 2.500 3.145 ;
        RECT  0.180 2.885 2.500 3.145 ;
        RECT  0.180 2.885 1.820 3.200 ;
        RECT  1.480 2.885 1.820 3.740 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  4.040 0.630 4.415 0.970 ;
        RECT  2.780 0.630 3.010 2.235 ;
        RECT  4.080 1.965 4.415 2.290 ;
        RECT  2.780 2.005 4.415 2.235 ;
        RECT  4.185 0.630 4.415 2.290 ;
        RECT  3.425 2.005 4.415 2.290 ;
        RECT  3.425 2.005 3.655 3.850 ;
        RECT  3.425 3.510 3.765 3.850 ;
        RECT  4.810 0.800 5.640 1.140 ;
        RECT  5.410 0.800 5.640 1.870 ;
        RECT  5.410 1.640 6.635 1.870 ;
        RECT  6.405 1.640 6.635 3.650 ;
        RECT  3.995 3.420 6.635 3.650 ;
        RECT  5.440 3.420 5.780 3.730 ;
        RECT  3.995 3.420 4.330 3.850 ;
        RECT  7.270 0.630 7.760 0.915 ;
        RECT  7.270 0.630 7.610 1.460 ;
        RECT  7.270 1.185 7.920 1.460 ;
        RECT  7.690 1.185 7.920 2.990 ;
        RECT  6.865 2.760 7.920 2.990 ;
        RECT  6.865 2.760 7.170 3.190 ;
        RECT  0.290 1.590 1.20 1.820 ;
        RECT  0.180 2.885 1.70 3.145 ;
        RECT  3.995 3.420 5.70 3.650 ;
    END
END NA7X0

MACRO NA6X4
    CLASS CORE ;
    FOREIGN NA6X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.975 0.505 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.470 2.030 4.220 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.265 2.120 8.735 2.640 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.793  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.215 1.125 7.695 1.465 ;
        RECT  7.215 1.125 7.570 3.930 ;
        RECT  5.790 2.550 7.570 2.780 ;
        RECT  7.055 2.250 7.570 2.780 ;
        RECT  5.915 1.240 6.255 2.780 ;
        RECT  5.790 2.550 6.130 3.930 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.985 1.620 9.325 2.830 ;
        RECT  8.945 1.620 9.325 2.025 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.075 3.470 10.585 4.250 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.430 3.580 9.770 5.280 ;
        RECT  7.950 3.090 8.290 5.280 ;
        RECT  6.510 3.010 6.850 5.280 ;
        RECT  4.560 2.560 5.370 5.280 ;
        RECT  2.260 2.560 2.600 5.280 ;
        RECT  0.740 4.095 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  8.075 -0.400 8.415 1.460 ;
        RECT  6.635 -0.400 6.975 1.550 ;
        RECT  5.055 -0.400 5.395 1.455 ;
        RECT  3.410 -0.400 3.790 1.575 ;
        RECT  1.840 -0.400 2.180 1.230 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.700 0.520 1.745 ;
        RECT  0.180 1.460 2.720 1.745 ;
        RECT  1.700 1.460 2.720 1.800 ;
        RECT  1.700 1.460 1.930 3.200 ;
        RECT  0.180 2.860 1.930 3.200 ;
        RECT  2.645 0.700 3.180 1.040 ;
        RECT  2.950 0.700 3.180 2.235 ;
        RECT  4.170 1.130 4.515 2.240 ;
        RECT  2.950 1.900 5.685 2.235 ;
        RECT  3.410 1.900 5.685 2.240 ;
        RECT  3.410 1.900 3.750 3.880 ;
        RECT  10.190 0.630 10.545 1.515 ;
        RECT  9.630 1.080 10.545 1.515 ;
        RECT  9.575 2.900 10.545 3.240 ;
        RECT  10.315 0.630 10.545 3.240 ;
        RECT  8.670 3.060 9.805 3.345 ;
        RECT  8.670 3.060 9.015 3.930 ;
        RECT  0.180 1.460 1.60 1.745 ;
        RECT  2.950 1.900 4.50 2.235 ;
        RECT  3.410 1.900 4.80 2.240 ;
    END
END NA6X4

MACRO NA6X2
    CLASS CORE ;
    FOREIGN NA6X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.975 0.505 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.340 3.470 2.030 4.065 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.755 2.130 6.220 2.630 ;
        RECT  5.755 2.120 6.215 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.815 1.640 5.545 2.020 ;
        RECT  4.815 1.260 5.175 2.020 ;
        RECT  4.815 1.260 5.170 3.700 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.560 1.620 6.920 2.145 ;
        RECT  6.425 1.620 6.920 2.025 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.555 3.470 8.065 4.130 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.870 3.600 7.210 5.280 ;
        RECT  5.550 2.860 5.890 5.280 ;
        RECT  4.110 2.780 4.450 5.280 ;
        RECT  2.260 2.780 2.600 5.280 ;
        RECT  0.740 3.595 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  5.630 -0.400 5.970 1.420 ;
        RECT  4.075 -0.400 4.415 1.670 ;
        RECT  3.410 -0.400 4.415 1.140 ;
        RECT  1.840 -0.400 2.180 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.350 2.720 1.690 ;
        RECT  1.700 1.350 2.720 1.800 ;
        RECT  1.700 1.350 1.930 3.200 ;
        RECT  0.180 2.860 1.930 3.200 ;
        RECT  2.645 0.700 3.180 1.040 ;
        RECT  2.950 0.700 3.180 2.235 ;
        RECT  2.950 1.900 3.970 2.235 ;
        RECT  3.410 1.900 3.970 2.240 ;
        RECT  3.410 1.900 3.750 4.100 ;
        RECT  7.670 0.630 8.025 1.470 ;
        RECT  7.670 0.630 7.900 3.200 ;
        RECT  6.310 2.860 8.015 3.200 ;
        RECT  0.180 1.350 1.20 1.690 ;
    END
END NA6X2

MACRO NA6X1
    CLASS CORE ;
    FOREIGN NA6X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.975 0.505 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.430 2.630 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.660 3.470 2.395 3.850 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.040 1.640 5.545 2.020 ;
        RECT  4.830 2.260 5.270 2.600 ;
        RECT  5.040 1.640 5.270 2.600 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 1.640 4.470 2.020 ;
        RECT  4.130 1.240 4.470 2.020 ;
        RECT  3.770 3.360 4.125 3.700 ;
        RECT  3.895 1.640 4.125 3.700 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.500 2.250 6.175 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.220 3.430 6.805 3.890 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.815 3.600 5.990 5.280 ;
        RECT  2.200 4.080 2.540 5.280 ;
        RECT  0.880 3.595 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.890 -0.400 5.230 0.960 ;
        RECT  3.395 -0.400 3.735 1.120 ;
        RECT  1.790 -0.400 2.130 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.350 2.650 1.690 ;
        RECT  0.290 2.860 1.890 3.090 ;
        RECT  1.660 1.350 1.890 3.200 ;
        RECT  1.440 2.860 1.890 3.200 ;
        RECT  0.290 2.860 0.520 3.940 ;
        RECT  0.180 3.600 0.520 3.940 ;
        RECT  2.595 0.780 3.110 1.120 ;
        RECT  2.880 0.780 3.110 2.490 ;
        RECT  2.880 2.260 3.665 2.490 ;
        RECT  3.190 2.260 3.665 2.600 ;
        RECT  3.190 2.260 3.530 3.120 ;
        RECT  6.410 1.360 6.750 1.700 ;
        RECT  6.410 1.360 6.640 3.200 ;
        RECT  5.090 2.860 6.755 3.200 ;
        RECT  4.355 2.970 6.755 3.200 ;
        RECT  2.950 3.820 3.290 4.160 ;
        RECT  4.355 2.970 4.585 4.160 ;
        RECT  2.950 3.930 4.585 4.160 ;
        RECT  0.180 1.350 1.30 1.690 ;
        RECT  4.355 2.970 5.20 3.200 ;
    END
END NA6X1

MACRO NA6X0
    CLASS CORE ;
    FOREIGN NA6X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.790 1.690 6.175 2.630 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.080 0.525 2.675 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.587  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.550 4.135 3.890 ;
        RECT  3.905 1.690 4.135 3.890 ;
        RECT  3.275 1.690 4.135 2.020 ;
        RECT  3.275 1.640 3.850 2.020 ;
        RECT  3.510 1.330 3.850 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 1.360 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 1.990 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.510 2.080 4.940 2.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.260 1.640 5.560 2.630 ;
        RECT  5.165 1.640 5.560 2.020 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.710 3.530 6.050 5.280 ;
        RECT  4.365 2.880 4.650 5.280 ;
        RECT  2.180 3.530 2.520 5.280 ;
        RECT  0.780 3.530 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.310 -0.400 4.650 1.470 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  2.220 1.260 2.500 3.165 ;
        RECT  0.180 2.905 2.500 3.165 ;
        RECT  0.180 2.905 1.820 3.220 ;
        RECT  1.480 2.905 1.820 3.760 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 3.870 ;
        RECT  3.360 2.250 3.675 2.590 ;
        RECT  2.780 2.360 3.675 2.590 ;
        RECT  2.780 2.360 3.045 3.870 ;
        RECT  2.780 3.530 3.335 3.870 ;
        RECT  6.295 0.630 6.690 1.470 ;
        RECT  6.310 2.880 6.690 3.220 ;
        RECT  6.405 0.630 6.690 3.220 ;
        RECT  5.010 2.935 6.690 3.220 ;
        RECT  5.010 2.935 5.350 3.760 ;
        RECT  0.290 1.590 1.50 1.820 ;
        RECT  0.180 2.905 1.10 3.165 ;
    END
END NA6X0

MACRO NA6I5X4
    CLASS CORE ;
    FOREIGN NA6I5X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.925 2.850 9.325 3.240 ;
        RECT  8.925 2.030 9.155 3.240 ;
        RECT  8.815 2.030 9.155 2.370 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.290 0.520 3.890 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.200 2.245 10.650 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.520 2.005 9.970 2.630 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 3.340 1.600 3.680 ;
        RECT  0.750 2.860 1.135 3.680 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.883  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.740 3.050 8.530 3.390 ;
        RECT  8.300 1.685 8.530 3.390 ;
        RECT  7.625 1.685 8.530 2.020 ;
        RECT  7.625 1.435 8.065 2.020 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.250 2.310 3.750 2.725 ;
        RECT  3.250 2.215 3.670 2.725 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.685 3.970 11.030 5.280 ;
        RECT  8.770 4.120 9.115 5.280 ;
        RECT  7.365 3.730 7.730 5.280 ;
        RECT  6.120 3.695 6.460 5.280 ;
        RECT  3.760 4.170 4.100 5.280 ;
        RECT  2.640 4.165 2.980 5.280 ;
        RECT  0.940 3.910 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.145 -0.400 10.970 0.855 ;
        RECT  8.385 -0.400 8.725 0.745 ;
        RECT  6.595 -0.400 6.935 1.180 ;
        RECT  4.790 -0.400 5.120 0.710 ;
        RECT  3.675 -0.400 4.015 0.710 ;
        RECT  0.880 -0.400 1.220 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.885 2.295 2.200 ;
        RECT  0.180 0.640 0.520 3.020 ;
        RECT  1.480 1.315 1.820 1.655 ;
        RECT  1.480 1.425 2.910 1.655 ;
        RECT  2.655 1.425 2.910 2.660 ;
        RECT  2.655 2.195 2.995 2.660 ;
        RECT  1.500 2.430 2.995 2.660 ;
        RECT  1.500 2.430 1.845 2.935 ;
        RECT  2.010 0.630 2.350 0.970 ;
        RECT  2.120 0.940 4.005 1.170 ;
        RECT  3.775 0.940 4.005 1.990 ;
        RECT  3.775 1.760 4.570 1.990 ;
        RECT  4.040 1.760 4.570 2.235 ;
        RECT  5.530 2.330 6.220 2.670 ;
        RECT  3.195 2.960 4.570 3.190 ;
        RECT  3.195 2.960 3.540 3.805 ;
        RECT  1.880 3.575 3.540 3.805 ;
        RECT  4.340 1.760 4.570 4.250 ;
        RECT  1.880 3.575 2.235 4.120 ;
        RECT  5.530 2.330 5.785 4.250 ;
        RECT  4.340 4.020 5.785 4.250 ;
        RECT  4.235 1.185 5.170 1.525 ;
        RECT  4.940 1.185 5.170 3.790 ;
        RECT  5.550 1.280 5.895 2.100 ;
        RECT  4.940 1.800 5.895 2.100 ;
        RECT  4.940 1.870 7.290 2.100 ;
        RECT  7.055 1.870 7.290 2.650 ;
        RECT  7.055 2.310 8.070 2.650 ;
        RECT  4.940 1.800 5.295 3.790 ;
        RECT  9.170 1.435 9.510 1.775 ;
        RECT  9.170 1.545 11.135 1.775 ;
        RECT  10.640 1.545 11.135 1.995 ;
        RECT  10.905 2.340 11.340 2.680 ;
        RECT  10.905 1.545 11.135 3.425 ;
        RECT  10.190 3.085 11.135 3.425 ;
        RECT  5.350 0.630 6.360 0.915 ;
        RECT  7.165 0.975 9.940 1.205 ;
        RECT  11.385 0.810 11.800 1.315 ;
        RECT  9.740 1.085 11.800 1.315 ;
        RECT  6.130 0.630 6.360 1.640 ;
        RECT  7.165 0.975 7.395 1.640 ;
        RECT  6.130 1.410 7.395 1.640 ;
        RECT  11.570 0.810 11.800 4.165 ;
        RECT  11.450 3.820 11.800 4.165 ;
        RECT  0.180 1.885 1.40 2.200 ;
        RECT  4.940 1.870 6.80 2.100 ;
        RECT  7.165 0.975 8.40 1.205 ;
        RECT  9.740 1.085 10.40 1.315 ;
    END
END NA6I5X4

MACRO NA6I5X2
    CLASS CORE ;
    FOREIGN NA6I5X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.885 7.435 3.240 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.250 0.760 3.850 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.310 2.245 8.760 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.885 8.080 2.630 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.395 3.340 1.775 3.835 ;
        RECT  1.260 3.340 1.775 3.805 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.575 1.640 6.805 3.395 ;
        RECT  6.275 3.160 6.615 4.080 ;
        RECT  6.410 1.640 6.805 2.020 ;
        RECT  6.060 1.640 6.805 1.870 ;
        RECT  6.060 1.110 6.400 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.370 1.620 3.715 2.700 ;
        RECT  3.265 1.620 3.715 2.035 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.795 3.970 9.140 5.280 ;
        RECT  7.035 4.085 7.380 5.280 ;
        RECT  5.550 3.730 5.905 5.280 ;
        RECT  3.695 3.700 4.035 5.280 ;
        RECT  2.115 2.955 2.780 3.300 ;
        RECT  2.005 3.810 2.350 5.280 ;
        RECT  2.115 2.955 2.350 5.280 ;
        RECT  0.940 4.035 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.580 -0.400 8.920 0.710 ;
        RECT  6.810 -0.400 7.155 0.970 ;
        RECT  5.270 -0.400 5.610 1.185 ;
        RECT  3.790 -0.400 4.130 0.710 ;
        RECT  0.915 -0.400 1.255 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.860 2.295 2.175 ;
        RECT  0.180 0.640 0.520 3.020 ;
        RECT  1.515 1.290 1.855 1.630 ;
        RECT  1.515 1.400 2.910 1.630 ;
        RECT  2.655 1.400 2.910 2.660 ;
        RECT  2.655 2.320 2.995 2.660 ;
        RECT  1.500 2.430 2.995 2.660 ;
        RECT  1.500 2.430 1.845 3.025 ;
        RECT  2.130 0.630 2.470 1.170 ;
        RECT  2.130 0.940 4.220 1.170 ;
        RECT  3.990 1.475 4.350 1.830 ;
        RECT  3.990 0.940 4.220 3.190 ;
        RECT  3.130 2.960 4.220 3.190 ;
        RECT  3.130 2.960 3.475 3.300 ;
        RECT  3.130 2.960 3.415 4.145 ;
        RECT  2.700 3.790 3.415 4.145 ;
        RECT  4.550 0.815 4.970 1.155 ;
        RECT  4.740 0.815 4.970 2.585 ;
        RECT  4.880 2.340 6.345 2.680 ;
        RECT  4.880 2.340 5.230 3.365 ;
        RECT  7.460 1.270 7.800 1.630 ;
        RECT  7.460 1.400 9.245 1.630 ;
        RECT  8.860 1.400 9.245 1.785 ;
        RECT  9.015 2.340 9.450 2.680 ;
        RECT  9.015 1.400 9.245 3.395 ;
        RECT  8.455 3.055 9.245 3.395 ;
        RECT  7.385 0.630 8.300 0.915 ;
        RECT  8.070 0.630 8.300 1.170 ;
        RECT  9.400 0.630 9.910 1.170 ;
        RECT  8.070 0.940 9.910 1.170 ;
        RECT  9.680 0.630 9.910 4.165 ;
        RECT  9.560 3.820 9.910 4.165 ;
        RECT  0.180 1.860 1.30 2.175 ;
        RECT  2.130 0.940 3.20 1.170 ;
    END
END NA6I5X2

MACRO NA6I5X1
    CLASS CORE ;
    FOREIGN NA6I5X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.920 6.805 3.240 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.250 0.760 3.850 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 2.245 8.130 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.885 7.450 2.630 ;
        END
    END BN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.395 3.340 1.825 3.835 ;
        RECT  1.315 3.340 1.825 3.800 ;
        RECT  1.260 3.340 1.825 3.680 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.781  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.945 1.640 6.175 3.165 ;
        RECT  5.645 2.930 5.985 3.800 ;
        RECT  5.780 1.640 6.175 2.020 ;
        RECT  5.370 1.640 6.175 1.870 ;
        RECT  5.370 1.480 5.710 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 1.495 3.850 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.155 3.970 8.500 5.280 ;
        RECT  6.405 4.085 6.750 5.280 ;
        RECT  4.115 3.900 4.455 5.280 ;
        RECT  2.795 3.730 3.135 5.280 ;
        RECT  0.940 4.035 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.685 -0.400 8.470 0.710 ;
        RECT  6.120 -0.400 6.460 0.970 ;
        RECT  5.390 -0.400 5.730 0.970 ;
        RECT  3.790 -0.400 4.130 0.710 ;
        RECT  0.915 -0.400 1.255 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.860 2.615 2.175 ;
        RECT  0.180 0.640 0.520 3.020 ;
        RECT  1.515 1.290 1.855 1.630 ;
        RECT  1.515 1.400 3.095 1.630 ;
        RECT  2.865 2.255 3.455 2.595 ;
        RECT  2.865 1.400 3.095 2.810 ;
        RECT  1.500 2.580 3.095 2.810 ;
        RECT  1.500 2.580 1.845 3.025 ;
        RECT  2.130 0.630 2.470 1.170 ;
        RECT  2.130 0.940 4.350 1.170 ;
        RECT  4.120 1.260 4.535 1.600 ;
        RECT  3.355 2.960 4.350 3.190 ;
        RECT  4.120 0.940 4.350 3.190 ;
        RECT  2.090 3.070 3.695 3.300 ;
        RECT  2.090 3.070 2.375 3.815 ;
        RECT  2.055 3.475 2.375 3.815 ;
        RECT  4.590 0.630 5.050 0.970 ;
        RECT  4.820 0.630 5.050 2.700 ;
        RECT  4.820 2.360 5.715 2.700 ;
        RECT  4.930 2.360 5.270 4.240 ;
        RECT  6.730 1.300 7.045 1.630 ;
        RECT  6.730 1.325 7.070 1.630 ;
        RECT  6.730 1.400 8.615 1.630 ;
        RECT  8.130 1.400 8.615 1.685 ;
        RECT  8.385 2.340 8.820 2.680 ;
        RECT  8.385 1.400 8.615 3.395 ;
        RECT  7.825 3.055 8.615 3.395 ;
        RECT  6.690 0.630 7.455 0.915 ;
        RECT  7.225 0.630 7.455 1.155 ;
        RECT  8.915 0.630 9.280 1.170 ;
        RECT  7.245 0.940 9.280 1.170 ;
        RECT  9.050 0.630 9.280 4.165 ;
        RECT  8.930 3.820 9.280 4.165 ;
        RECT  0.180 1.860 1.50 2.175 ;
        RECT  2.130 0.940 3.00 1.170 ;
        RECT  7.245 0.940 8.40 1.170 ;
    END
END NA6I5X1

MACRO NA6I5X0
    CLASS CORE ;
    FOREIGN NA6I5X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.210 0.800 3.550 ;
        RECT  0.125 3.210 0.505 3.965 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 2.240 8.115 2.790 ;
        END
    END AN
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.405 3.340 1.825 3.820 ;
        RECT  1.300 3.340 1.825 3.800 ;
        END
    END EN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.585  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.750 3.620 6.175 3.960 ;
        RECT  5.945 1.640 6.175 3.960 ;
        RECT  5.280 1.640 6.175 2.020 ;
        RECT  5.280 1.365 5.620 2.020 ;
        END
    END Q
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.405 2.860 6.805 3.240 ;
        RECT  6.405 1.980 6.740 3.240 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.860 7.440 2.630 ;
        END
    END BN
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 1.495 3.840 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.815 3.530 9.155 5.280 ;
        RECT  6.450 3.575 6.790 5.280 ;
        RECT  4.220 3.530 4.560 5.280 ;
        RECT  2.820 3.530 3.160 5.280 ;
        RECT  0.980 4.035 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.645 -0.400 8.465 0.710 ;
        RECT  6.080 -0.400 6.420 0.970 ;
        RECT  5.380 -0.400 5.720 0.970 ;
        RECT  3.780 -0.400 4.120 0.710 ;
        RECT  0.880 -0.400 1.220 0.870 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.860 2.635 2.175 ;
        RECT  0.180 0.630 0.520 2.980 ;
        RECT  1.480 1.170 1.820 1.630 ;
        RECT  1.480 1.400 3.095 1.630 ;
        RECT  2.865 2.250 3.610 2.540 ;
        RECT  2.865 1.400 3.095 2.810 ;
        RECT  1.645 2.525 3.095 2.810 ;
        RECT  1.645 2.525 1.985 2.925 ;
        RECT  2.120 0.630 2.460 1.170 ;
        RECT  2.120 0.940 4.350 1.170 ;
        RECT  4.120 0.940 4.350 1.490 ;
        RECT  2.165 3.070 4.590 3.300 ;
        RECT  4.300 1.260 4.590 3.300 ;
        RECT  2.130 3.105 2.360 3.850 ;
        RECT  3.520 3.070 3.860 3.760 ;
        RECT  2.055 3.510 2.360 3.850 ;
        RECT  4.580 0.630 5.050 0.970 ;
        RECT  4.820 0.630 5.050 2.700 ;
        RECT  4.820 2.360 5.715 2.700 ;
        RECT  5.035 2.360 5.375 3.870 ;
        RECT  6.680 1.300 6.995 1.610 ;
        RECT  6.680 1.270 6.965 1.610 ;
        RECT  6.735 1.400 8.615 1.630 ;
        RECT  8.080 1.400 8.615 1.685 ;
        RECT  8.385 1.865 8.820 2.205 ;
        RECT  8.385 1.400 8.615 3.400 ;
        RECT  8.010 3.115 8.615 3.400 ;
        RECT  8.010 3.115 8.350 3.455 ;
        RECT  6.690 0.630 7.415 0.915 ;
        RECT  7.185 0.630 7.415 1.170 ;
        RECT  7.185 0.940 9.280 1.170 ;
        RECT  8.925 0.940 9.280 1.280 ;
        RECT  9.050 0.940 9.280 3.070 ;
        RECT  8.845 2.730 9.280 3.070 ;
        RECT  0.180 1.860 1.80 2.175 ;
        RECT  2.120 0.940 3.40 1.170 ;
        RECT  2.165 3.070 3.90 3.300 ;
        RECT  7.185 0.940 8.40 1.170 ;
    END
END NA6I5X0

MACRO NA6I4X4
    CLASS CORE ;
    FOREIGN NA6I4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.295 2.850 8.695 3.240 ;
        RECT  8.295 2.030 8.525 3.240 ;
        RECT  8.185 2.030 8.525 2.370 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.070 0.675 2.410 ;
        RECT  0.120 2.070 0.530 3.250 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.570 2.245 10.020 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.890 2.005 9.340 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.883  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.110 3.050 7.900 3.390 ;
        RECT  7.670 1.685 7.900 3.390 ;
        RECT  6.995 1.685 7.900 2.020 ;
        RECT  6.995 1.435 7.435 2.020 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.305 3.125 2.730 ;
        RECT  2.635 2.210 3.045 2.730 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 1.625 2.405 2.540 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.055 3.970 10.400 5.280 ;
        RECT  8.140 4.120 8.485 5.280 ;
        RECT  6.735 3.730 7.100 5.280 ;
        RECT  5.490 3.695 5.830 5.280 ;
        RECT  3.130 4.170 3.470 5.280 ;
        RECT  2.010 4.165 2.350 5.280 ;
        RECT  0.230 3.480 0.570 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  9.515 -0.400 10.340 0.855 ;
        RECT  7.755 -0.400 8.095 0.745 ;
        RECT  5.965 -0.400 6.305 1.180 ;
        RECT  4.160 -0.400 4.490 0.710 ;
        RECT  3.045 -0.400 3.385 0.710 ;
        RECT  0.250 -0.400 0.590 1.005 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.850 1.315 1.190 1.655 ;
        RECT  0.960 2.080 1.745 2.425 ;
        RECT  0.960 1.315 1.190 2.980 ;
        RECT  0.790 2.640 1.190 2.980 ;
        RECT  1.380 0.630 1.720 0.970 ;
        RECT  1.490 0.940 3.375 1.170 ;
        RECT  3.145 0.940 3.375 1.990 ;
        RECT  3.145 1.760 3.940 1.990 ;
        RECT  3.410 1.760 3.940 2.235 ;
        RECT  4.900 2.330 5.590 2.670 ;
        RECT  2.565 2.960 3.940 3.190 ;
        RECT  2.565 2.960 2.910 3.600 ;
        RECT  1.250 3.370 2.910 3.600 ;
        RECT  2.570 2.960 2.910 3.770 ;
        RECT  3.710 1.760 3.940 4.250 ;
        RECT  1.250 3.370 1.605 4.180 ;
        RECT  4.900 2.330 5.155 4.250 ;
        RECT  3.710 4.020 5.155 4.250 ;
        RECT  3.605 1.185 4.540 1.525 ;
        RECT  4.310 1.185 4.540 3.790 ;
        RECT  4.920 1.280 5.265 2.100 ;
        RECT  4.310 1.800 5.265 2.100 ;
        RECT  4.310 1.870 6.660 2.100 ;
        RECT  6.425 1.870 6.660 2.650 ;
        RECT  6.425 2.310 7.440 2.650 ;
        RECT  4.310 1.800 4.665 3.790 ;
        RECT  8.540 1.435 8.880 1.775 ;
        RECT  8.540 1.545 10.505 1.775 ;
        RECT  10.010 1.545 10.505 1.995 ;
        RECT  10.275 2.340 10.710 2.680 ;
        RECT  10.275 1.545 10.505 3.425 ;
        RECT  9.560 3.085 10.505 3.425 ;
        RECT  4.720 0.630 5.730 0.915 ;
        RECT  6.535 0.975 9.310 1.205 ;
        RECT  10.755 0.810 11.170 1.315 ;
        RECT  9.110 1.085 11.170 1.315 ;
        RECT  5.500 0.630 5.730 1.640 ;
        RECT  6.535 0.975 6.765 1.640 ;
        RECT  5.500 1.410 6.765 1.640 ;
        RECT  10.940 0.810 11.170 4.165 ;
        RECT  10.820 3.820 11.170 4.165 ;
        RECT  4.310 1.870 5.90 2.100 ;
        RECT  6.535 0.975 8.30 1.205 ;
        RECT  9.110 1.085 10.20 1.315 ;
    END
END NA6I4X4

MACRO NA6I4X2
    CLASS CORE ;
    FOREIGN NA6I4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.885 6.805 3.240 ;
        END
    END CN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 2.245 8.130 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.885 7.450 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.945 1.640 6.175 3.395 ;
        RECT  5.645 3.160 5.985 4.080 ;
        RECT  5.780 1.640 6.175 2.020 ;
        RECT  5.430 1.640 6.175 1.870 ;
        RECT  5.430 1.110 5.770 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.740 1.620 3.085 2.700 ;
        RECT  2.635 1.620 3.085 2.035 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.940 2.195 2.460 2.675 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.640 2.640 ;
        END
    END DN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.165 3.970 8.510 5.280 ;
        RECT  6.405 4.085 6.750 5.280 ;
        RECT  4.920 3.730 5.275 5.280 ;
        RECT  3.065 3.700 3.405 5.280 ;
        RECT  1.485 2.955 2.150 3.300 ;
        RECT  1.355 3.810 1.720 5.280 ;
        RECT  1.485 2.955 1.720 5.280 ;
        RECT  0.310 3.455 0.650 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.950 -0.400 8.290 0.710 ;
        RECT  6.180 -0.400 6.525 0.970 ;
        RECT  4.640 -0.400 4.980 1.185 ;
        RECT  3.160 -0.400 3.500 0.710 ;
        RECT  0.285 -0.400 0.625 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.870 1.290 1.230 2.175 ;
        RECT  0.870 1.835 1.665 2.175 ;
        RECT  0.870 1.290 1.215 3.025 ;
        RECT  1.500 0.630 1.840 1.170 ;
        RECT  1.500 0.940 3.720 1.170 ;
        RECT  3.360 1.475 3.720 1.830 ;
        RECT  3.490 0.940 3.720 3.190 ;
        RECT  2.500 2.960 3.720 3.190 ;
        RECT  2.500 2.960 2.845 3.300 ;
        RECT  2.500 2.960 2.785 4.145 ;
        RECT  2.070 3.790 2.785 4.145 ;
        RECT  3.950 0.720 4.340 1.060 ;
        RECT  4.110 0.720 4.340 2.585 ;
        RECT  4.250 2.340 5.715 2.680 ;
        RECT  4.250 2.340 4.600 3.365 ;
        RECT  6.830 1.270 7.170 1.630 ;
        RECT  6.830 1.400 8.615 1.630 ;
        RECT  8.230 1.400 8.615 1.785 ;
        RECT  8.385 2.340 8.820 2.680 ;
        RECT  8.385 1.400 8.615 3.395 ;
        RECT  7.825 3.055 8.615 3.395 ;
        RECT  6.755 0.630 7.670 0.915 ;
        RECT  7.440 0.630 7.670 1.170 ;
        RECT  8.770 0.630 9.280 1.170 ;
        RECT  7.440 0.940 9.280 1.170 ;
        RECT  9.050 0.630 9.280 4.135 ;
        RECT  8.930 3.790 9.280 4.135 ;
        RECT  1.500 0.940 2.80 1.170 ;
    END
END NA6I4X2

MACRO NA6I4X1
    CLASS CORE ;
    FOREIGN NA6I4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 2.250 2.195 2.630 ;
        END
    END E
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.920 5.545 3.240 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.560 2.210 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.420 2.240 6.870 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.885 6.190 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.685 1.640 4.915 3.165 ;
        RECT  4.385 2.930 4.725 3.805 ;
        RECT  4.525 1.640 4.915 2.020 ;
        RECT  4.110 1.640 4.915 1.875 ;
        RECT  4.110 1.480 4.450 1.875 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.495 2.590 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.895 3.970 7.240 5.280 ;
        RECT  5.145 4.085 5.490 5.280 ;
        RECT  2.855 3.900 3.195 5.280 ;
        RECT  0.900 3.790 1.710 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.425 -0.400 7.210 0.710 ;
        RECT  4.860 -0.400 5.200 0.970 ;
        RECT  4.130 -0.400 4.470 0.970 ;
        RECT  2.530 -0.400 2.870 0.710 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.790 1.425 1.120 2.460 ;
        RECT  0.790 2.110 1.205 2.460 ;
        RECT  0.290 2.440 1.065 2.670 ;
        RECT  0.290 2.440 0.520 4.125 ;
        RECT  0.180 3.785 0.520 4.125 ;
        RECT  0.910 0.720 1.250 1.170 ;
        RECT  0.910 0.940 3.090 1.170 ;
        RECT  2.860 1.260 3.275 1.600 ;
        RECT  0.775 2.905 1.120 3.300 ;
        RECT  2.095 2.960 3.090 3.190 ;
        RECT  2.860 0.940 3.090 3.190 ;
        RECT  0.775 3.070 2.435 3.300 ;
        RECT  3.330 0.630 3.790 0.970 ;
        RECT  3.560 0.630 3.790 2.700 ;
        RECT  3.560 2.360 4.455 2.700 ;
        RECT  3.670 2.360 3.935 4.240 ;
        RECT  3.670 3.900 4.010 4.240 ;
        RECT  5.470 1.300 5.785 1.630 ;
        RECT  5.470 1.325 5.810 1.630 ;
        RECT  5.470 1.400 7.355 1.630 ;
        RECT  6.870 1.400 7.355 1.685 ;
        RECT  7.125 2.340 7.560 2.680 ;
        RECT  7.125 1.400 7.355 3.395 ;
        RECT  6.565 3.055 7.355 3.395 ;
        RECT  5.430 0.630 6.195 0.915 ;
        RECT  5.965 0.630 6.195 1.155 ;
        RECT  7.655 0.630 8.020 1.170 ;
        RECT  5.985 0.940 8.020 1.170 ;
        RECT  7.790 0.630 8.020 4.165 ;
        RECT  7.670 3.820 8.020 4.165 ;
        RECT  0.910 0.940 2.60 1.170 ;
        RECT  5.985 0.940 7.30 1.170 ;
    END
END NA6I4X1

MACRO NA6I4X0
    CLASS CORE ;
    FOREIGN NA6I4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.915 0.605 2.630 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.593  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.490 3.620 4.915 3.960 ;
        RECT  4.685 1.640 4.915 3.960 ;
        RECT  4.020 1.640 4.915 2.020 ;
        RECT  4.020 1.330 4.360 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.785 0.945 2.395 1.360 ;
        RECT  1.785 0.630 2.125 1.360 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.360 2.050 3.025 2.630 ;
        END
    END F
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 2.860 5.545 3.240 ;
        RECT  5.145 1.975 5.480 3.240 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.860 6.180 2.630 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 2.235 6.845 2.795 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.555 3.530 7.895 5.280 ;
        RECT  5.190 3.770 5.530 5.280 ;
        RECT  2.960 3.530 3.300 5.280 ;
        RECT  1.560 3.960 1.900 5.280 ;
        RECT  0.180 3.315 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.375 -0.400 7.205 0.710 ;
        RECT  4.820 -0.400 5.160 0.970 ;
        RECT  4.040 -0.400 4.380 0.970 ;
        RECT  2.440 -0.400 2.780 0.710 ;
        RECT  0.190 -0.400 0.530 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.195 1.170 0.535 1.510 ;
        RECT  0.195 1.225 1.065 1.510 ;
        RECT  0.835 1.225 1.065 2.980 ;
        RECT  0.835 2.050 1.600 2.335 ;
        RECT  0.835 2.050 1.120 2.980 ;
        RECT  1.120 0.630 1.555 0.970 ;
        RECT  1.325 0.630 1.555 1.820 ;
        RECT  3.040 1.155 3.330 1.820 ;
        RECT  1.325 1.590 3.330 1.820 ;
        RECT  1.830 1.590 2.060 3.440 ;
        RECT  0.940 3.210 2.600 3.440 ;
        RECT  0.940 3.210 1.280 3.680 ;
        RECT  2.260 3.210 2.600 3.760 ;
        RECT  3.240 0.630 3.790 0.925 ;
        RECT  3.560 0.630 3.790 2.700 ;
        RECT  3.560 2.360 4.455 2.700 ;
        RECT  3.775 2.360 4.115 3.870 ;
        RECT  5.420 1.300 5.725 1.610 ;
        RECT  5.420 1.270 5.705 1.610 ;
        RECT  5.475 1.400 7.305 1.630 ;
        RECT  6.820 1.400 7.305 1.685 ;
        RECT  7.075 1.865 7.560 2.205 ;
        RECT  7.075 1.400 7.305 3.455 ;
        RECT  6.750 3.115 7.305 3.455 ;
        RECT  5.560 0.630 6.145 0.915 ;
        RECT  5.915 0.630 6.145 1.170 ;
        RECT  5.915 0.940 8.020 1.170 ;
        RECT  7.665 0.940 8.020 1.280 ;
        RECT  7.790 0.940 8.020 3.070 ;
        RECT  7.555 2.730 8.020 3.070 ;
        RECT  1.325 1.590 2.20 1.820 ;
        RECT  5.915 0.940 7.50 1.170 ;
    END
END NA6I4X0

MACRO NA6I3X4
    CLASS CORE ;
    FOREIGN NA6I3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.310 2.245 8.860 3.070 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.625 2.090 8.080 2.635 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.986  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.480 2.970 6.820 4.180 ;
        RECT  6.410 1.530 6.815 2.030 ;
        RECT  6.410 1.530 6.640 3.390 ;
        RECT  5.120 3.050 6.820 3.390 ;
        RECT  5.895 1.530 6.815 1.780 ;
        RECT  5.895 1.435 6.235 1.780 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.230 2.035 2.710 ;
        END
    END F
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.850 7.435 3.240 ;
        RECT  7.055 2.310 7.285 3.240 ;
        RECT  6.925 2.310 7.285 2.650 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.700 0.550 3.270 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 1.625 1.145 2.520 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.795 3.955 9.140 5.280 ;
        RECT  5.715 3.730 6.080 5.280 ;
        RECT  4.400 3.045 4.740 5.280 ;
        RECT  2.060 4.170 2.400 5.280 ;
        RECT  0.940 4.165 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.255 -0.400 9.080 0.855 ;
        RECT  6.655 -0.400 6.995 0.745 ;
        RECT  4.865 -0.400 5.205 1.180 ;
        RECT  3.085 -0.400 3.415 0.710 ;
        RECT  1.970 -0.400 2.310 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.340 0.965 0.680 1.395 ;
        RECT  0.340 1.165 2.115 1.395 ;
        RECT  1.885 1.165 2.115 1.990 ;
        RECT  1.885 1.760 2.925 1.990 ;
        RECT  2.335 1.760 2.925 2.235 ;
        RECT  3.900 2.330 4.500 2.665 ;
        RECT  1.495 2.960 2.925 3.190 ;
        RECT  1.495 2.960 1.840 3.770 ;
        RECT  0.180 3.540 1.840 3.770 ;
        RECT  0.180 3.540 0.535 3.900 ;
        RECT  2.695 1.760 2.925 4.250 ;
        RECT  3.900 2.330 4.155 4.250 ;
        RECT  2.695 4.020 4.155 4.250 ;
        RECT  2.530 1.185 3.470 1.525 ;
        RECT  3.240 1.185 3.470 3.790 ;
        RECT  3.850 1.280 4.175 2.100 ;
        RECT  3.240 1.830 4.175 2.100 ;
        RECT  3.240 1.870 5.400 2.100 ;
        RECT  5.165 1.870 5.400 2.650 ;
        RECT  5.165 2.310 6.180 2.650 ;
        RECT  3.240 1.830 3.595 3.790 ;
        RECT  7.280 1.435 7.620 1.775 ;
        RECT  7.280 1.545 9.340 1.775 ;
        RECT  8.750 1.545 9.340 1.995 ;
        RECT  9.110 2.200 9.505 2.540 ;
        RECT  9.110 1.545 9.340 3.725 ;
        RECT  7.180 3.470 9.340 3.725 ;
        RECT  7.180 3.470 7.545 3.810 ;
        RECT  3.645 0.630 4.635 0.950 ;
        RECT  5.435 0.975 8.050 1.205 ;
        RECT  9.495 0.810 9.965 1.315 ;
        RECT  7.850 1.085 9.965 1.315 ;
        RECT  4.405 0.630 4.635 1.640 ;
        RECT  5.435 0.975 5.665 1.640 ;
        RECT  4.405 1.410 5.665 1.640 ;
        RECT  9.570 3.240 9.965 4.165 ;
        RECT  9.735 0.810 9.965 4.165 ;
        RECT  9.560 3.800 9.965 4.165 ;
        RECT  3.240 1.870 4.00 2.100 ;
        RECT  7.280 1.545 8.40 1.775 ;
        RECT  7.180 3.470 8.60 3.725 ;
        RECT  5.435 0.975 7.50 1.205 ;
        RECT  7.850 1.085 8.10 1.315 ;
    END
END NA6I3X4

MACRO NA6I3X2
    CLASS CORE ;
    FOREIGN NA6I3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.885 5.545 3.240 ;
        END
    END CN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.420 2.245 6.870 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.885 6.190 2.630 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.425 0.680 1.790 ;
        RECT  0.115 1.425 0.535 2.030 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.685 1.640 4.915 3.395 ;
        RECT  4.385 3.160 4.725 4.080 ;
        RECT  4.520 1.640 4.915 2.020 ;
        RECT  4.170 1.640 4.915 1.870 ;
        RECT  4.170 1.110 4.510 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.570 2.285 1.910 2.625 ;
        RECT  1.570 1.620 1.870 2.625 ;
        RECT  1.375 1.620 1.870 2.035 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 2.200 1.210 2.650 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.905 3.970 7.250 5.280 ;
        RECT  5.145 4.085 5.490 5.280 ;
        RECT  3.660 3.730 4.015 5.280 ;
        RECT  1.890 3.625 2.230 5.280 ;
        RECT  0.180 2.880 0.975 3.225 ;
        RECT  0.180 2.880 0.545 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.690 -0.400 7.030 0.710 ;
        RECT  4.920 -0.400 5.265 0.970 ;
        RECT  3.380 -0.400 3.720 1.185 ;
        RECT  1.900 -0.400 2.240 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.830 0.620 1.170 ;
        RECT  0.280 0.940 2.460 1.170 ;
        RECT  2.100 1.475 2.460 1.830 ;
        RECT  2.230 0.940 2.460 3.225 ;
        RECT  1.240 2.885 2.460 3.225 ;
        RECT  1.240 2.885 1.525 4.145 ;
        RECT  0.895 3.790 1.525 4.145 ;
        RECT  2.690 0.720 3.080 1.060 ;
        RECT  2.850 0.720 3.080 2.585 ;
        RECT  3.075 2.340 4.455 2.680 ;
        RECT  3.075 2.340 3.425 3.365 ;
        RECT  5.570 1.270 5.910 1.630 ;
        RECT  5.570 1.400 7.355 1.630 ;
        RECT  6.970 1.400 7.355 1.785 ;
        RECT  7.125 2.340 7.560 2.680 ;
        RECT  7.125 1.400 7.355 3.395 ;
        RECT  6.565 3.055 7.355 3.395 ;
        RECT  5.495 0.630 6.410 0.915 ;
        RECT  6.180 0.630 6.410 1.170 ;
        RECT  7.510 0.630 8.020 1.170 ;
        RECT  6.180 0.940 8.020 1.170 ;
        RECT  7.790 0.630 8.020 4.135 ;
        RECT  7.670 3.790 8.020 4.135 ;
        RECT  0.280 0.940 1.40 1.170 ;
    END
END NA6I3X2

MACRO NA6I3X1
    CLASS CORE ;
    FOREIGN NA6I3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.505 0.630 2.020 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.920 4.915 3.240 ;
        END
    END CN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.790 2.245 6.240 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.885 5.560 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.165 ;
        RECT  3.755 2.930 4.100 3.800 ;
        RECT  3.475 1.640 4.285 2.020 ;
        RECT  3.475 1.480 3.820 2.020 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.495 1.960 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.265 3.970 6.610 5.280 ;
        RECT  4.515 4.085 4.860 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.740 3.700 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.795 -0.400 6.580 0.710 ;
        RECT  4.230 -0.400 4.570 0.970 ;
        RECT  3.500 -0.400 3.840 0.970 ;
        RECT  1.900 -0.400 2.240 0.765 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.885 0.625 1.225 ;
        RECT  0.280 0.995 2.460 1.225 ;
        RECT  2.230 1.260 2.645 1.600 ;
        RECT  2.230 0.995 2.460 3.155 ;
        RECT  0.180 2.925 2.460 3.155 ;
        RECT  0.180 2.925 1.845 3.265 ;
        RECT  1.505 2.925 1.845 4.040 ;
        RECT  2.700 0.630 3.160 0.970 ;
        RECT  2.930 0.630 3.160 4.240 ;
        RECT  2.930 2.360 3.825 2.700 ;
        RECT  2.930 2.360 3.195 4.240 ;
        RECT  2.930 3.900 3.380 4.240 ;
        RECT  4.840 1.300 5.155 1.630 ;
        RECT  4.840 1.325 5.180 1.630 ;
        RECT  4.840 1.400 6.725 1.630 ;
        RECT  6.240 1.400 6.725 1.685 ;
        RECT  6.495 2.340 6.930 2.680 ;
        RECT  6.495 1.400 6.725 3.395 ;
        RECT  5.935 3.055 6.725 3.395 ;
        RECT  4.800 0.630 5.565 0.915 ;
        RECT  5.335 0.630 5.565 1.155 ;
        RECT  7.025 0.630 7.390 1.170 ;
        RECT  5.355 0.940 7.390 1.170 ;
        RECT  7.160 0.630 7.390 4.165 ;
        RECT  7.040 3.820 7.390 4.165 ;
        RECT  0.280 0.995 1.60 1.225 ;
        RECT  0.180 2.925 1.40 3.155 ;
        RECT  5.355 0.940 6.80 1.170 ;
    END
END NA6I3X1

MACRO NA6I3X0
    CLASS CORE ;
    FOREIGN NA6I3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.725 2.245 6.180 2.790 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.505 2.675 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.591  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.620 4.105 3.960 ;
        RECT  3.875 1.740 4.105 3.960 ;
        RECT  3.240 1.740 4.105 2.020 ;
        RECT  3.240 1.330 3.655 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 1.360 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 1.990 2.630 ;
        END
    END F
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.360 2.860 4.915 3.240 ;
        RECT  4.360 1.975 4.700 3.240 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.090 1.860 5.495 2.630 ;
        END
    END BN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.035 -0.400 7.375 0.710 ;
        RECT  5.600 -0.400 5.940 0.710 ;
        RECT  4.040 -0.400 4.380 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.985 3.440 7.325 5.280 ;
        RECT  4.410 3.770 4.750 5.280 ;
        RECT  2.180 3.530 2.520 5.280 ;
        RECT  0.780 3.515 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  0.735 1.590 0.965 3.220 ;
        RECT  0.180 2.905 0.965 3.220 ;
        RECT  0.180 2.935 1.710 3.220 ;
        RECT  1.480 2.935 1.710 3.760 ;
        RECT  1.480 3.420 1.820 3.760 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 3.870 ;
        RECT  2.780 2.360 3.645 2.700 ;
        RECT  2.780 2.360 3.045 3.870 ;
        RECT  2.780 3.530 3.335 3.870 ;
        RECT  4.640 1.300 4.950 1.610 ;
        RECT  4.640 1.270 4.925 1.610 ;
        RECT  4.695 1.400 6.755 1.630 ;
        RECT  6.040 1.400 6.755 1.685 ;
        RECT  6.515 1.855 6.830 2.195 ;
        RECT  6.515 1.400 6.755 3.455 ;
        RECT  5.970 3.115 6.755 3.455 ;
        RECT  4.650 0.630 5.370 0.915 ;
        RECT  5.140 0.630 5.370 1.170 ;
        RECT  5.140 0.940 7.290 1.170 ;
        RECT  7.035 1.170 7.375 1.510 ;
        RECT  7.060 1.170 7.375 2.990 ;
        RECT  7.005 2.640 7.375 2.990 ;
        RECT  0.290 1.590 1.40 1.820 ;
        RECT  4.695 1.400 5.40 1.630 ;
        RECT  5.140 0.940 6.30 1.170 ;
    END
END NA6I3X0

MACRO NA6I2X4
    CLASS CORE ;
    FOREIGN NA6I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.565 1.590 10.115 1.985 ;
        RECT  9.565 1.590 9.995 2.055 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.881  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.025 3.050 6.825 3.390 ;
        RECT  6.595 1.630 6.825 3.390 ;
        RECT  6.025 1.630 6.825 2.020 ;
        RECT  6.025 1.435 6.370 2.020 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 2.230 2.090 2.710 ;
        END
    END F
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.185 2.240 10.735 2.630 ;
        RECT  10.395 2.075 10.735 2.630 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.220 0.520 3.000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.205 2.540 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.875 7.445 3.240 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.100 2.860 10.440 5.280 ;
        RECT  8.175 4.170 8.515 5.280 ;
        RECT  7.055 4.170 7.400 5.280 ;
        RECT  5.650 3.730 6.015 5.280 ;
        RECT  4.405 3.695 4.745 5.280 ;
        RECT  0.945 4.165 2.405 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.015 -0.400 10.370 1.360 ;
        RECT  6.785 -0.400 7.125 0.710 ;
        RECT  4.995 -0.400 5.335 1.180 ;
        RECT  3.165 -0.400 3.495 0.710 ;
        RECT  1.980 -0.400 2.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.310 0.630 0.650 1.420 ;
        RECT  0.310 1.180 2.310 1.410 ;
        RECT  0.310 1.180 0.655 1.420 ;
        RECT  0.310 0.630 0.640 1.430 ;
        RECT  2.080 1.180 2.310 1.990 ;
        RECT  2.080 1.760 2.875 1.990 ;
        RECT  2.415 1.760 2.875 2.235 ;
        RECT  3.920 2.330 4.505 2.670 ;
        RECT  1.500 2.960 2.875 3.190 ;
        RECT  1.500 2.960 1.845 3.600 ;
        RECT  0.180 3.370 1.845 3.600 ;
        RECT  1.505 2.960 1.845 3.770 ;
        RECT  2.645 1.760 2.875 4.250 ;
        RECT  0.180 3.370 0.535 4.180 ;
        RECT  3.920 2.330 4.175 4.250 ;
        RECT  2.645 4.020 4.175 4.250 ;
        RECT  2.610 1.185 3.495 1.525 ;
        RECT  3.255 1.185 3.495 3.790 ;
        RECT  3.925 1.280 4.270 2.100 ;
        RECT  3.255 1.800 4.270 2.100 ;
        RECT  3.255 1.870 5.595 2.100 ;
        RECT  5.360 1.870 5.595 2.650 ;
        RECT  5.360 2.310 6.365 2.650 ;
        RECT  3.255 1.800 3.595 3.790 ;
        RECT  3.725 0.630 4.735 0.950 ;
        RECT  5.565 0.975 8.835 1.205 ;
        RECT  4.505 0.630 4.735 1.640 ;
        RECT  8.495 0.720 8.835 1.590 ;
        RECT  5.565 0.975 5.795 1.640 ;
        RECT  4.505 1.410 5.795 1.640 ;
        RECT  7.685 0.975 7.915 3.760 ;
        RECT  7.615 3.420 9.275 3.760 ;
        RECT  9.105 1.020 9.555 1.360 ;
        RECT  8.145 2.200 9.335 2.540 ;
        RECT  9.105 1.020 9.335 2.935 ;
        RECT  9.105 2.585 9.685 2.935 ;
        RECT  10.810 1.020 11.225 1.370 ;
        RECT  10.995 1.020 11.225 3.215 ;
        RECT  10.820 2.860 11.050 4.110 ;
        RECT  10.670 3.765 11.050 4.110 ;
        RECT  0.310 1.180 1.20 1.410 ;
        RECT  3.255 1.870 4.80 2.100 ;
        RECT  5.565 0.975 7.80 1.205 ;
    END
END NA6I2X4

MACRO NA6I2X2
    CLASS CORE ;
    FOREIGN NA6I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.530 0.630 2.020 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.635 1.575 8.170 2.045 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.270 2.805 8.795 3.285 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.955 5.510 3.240 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.685 1.640 4.915 3.360 ;
        RECT  4.475 3.125 4.815 4.045 ;
        RECT  4.535 1.640 4.915 2.020 ;
        RECT  4.270 1.150 4.610 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.575 1.960 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.210 3.680 8.550 5.280 ;
        RECT  6.360 3.705 6.700 5.280 ;
        RECT  5.235 3.705 5.580 5.280 ;
        RECT  3.715 4.065 4.055 5.280 ;
        RECT  0.885 3.635 2.345 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.115 -0.400 8.470 1.150 ;
        RECT  5.020 -0.400 5.370 1.035 ;
        RECT  3.500 -0.400 3.840 1.220 ;
        RECT  1.900 -0.400 2.240 0.785 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.960 0.620 1.300 ;
        RECT  0.280 1.070 2.460 1.300 ;
        RECT  2.230 1.480 2.660 1.825 ;
        RECT  2.230 1.070 2.460 3.090 ;
        RECT  0.180 2.860 2.460 3.090 ;
        RECT  1.445 2.860 1.785 3.235 ;
        RECT  0.180 2.860 0.520 3.985 ;
        RECT  2.700 0.720 3.160 1.060 ;
        RECT  2.930 0.720 3.160 2.700 ;
        RECT  2.930 2.455 4.455 2.700 ;
        RECT  3.200 2.455 4.455 2.795 ;
        RECT  3.200 2.455 3.540 3.675 ;
        RECT  5.600 0.630 5.985 0.915 ;
        RECT  5.740 0.630 5.985 1.775 ;
        RECT  5.740 1.435 7.145 1.775 ;
        RECT  5.740 0.630 5.970 3.290 ;
        RECT  7.130 2.880 7.470 3.290 ;
        RECT  5.740 2.950 7.470 3.290 ;
        RECT  6.565 0.720 7.690 1.060 ;
        RECT  6.930 3.535 7.830 3.875 ;
        RECT  7.490 3.535 7.830 4.040 ;
        RECT  8.930 0.810 9.270 1.150 ;
        RECT  6.200 2.330 9.270 2.565 ;
        RECT  6.200 2.330 6.490 2.700 ;
        RECT  9.040 0.810 9.270 4.040 ;
        RECT  8.930 3.695 9.270 4.040 ;
        RECT  0.280 1.070 1.80 1.300 ;
        RECT  0.180 2.860 1.30 3.090 ;
        RECT  6.200 2.330 8.70 2.565 ;
    END
END NA6I2X2

MACRO NA6I2X1
    CLASS CORE ;
    FOREIGN NA6I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.505 0.630 2.020 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.005 1.575 7.540 2.045 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.640 2.805 8.165 3.285 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.955 4.865 3.240 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.165 ;
        RECT  3.755 2.930 4.095 3.800 ;
        RECT  3.905 1.640 4.285 2.020 ;
        RECT  3.480 1.640 4.285 1.870 ;
        RECT  3.480 1.480 3.820 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.495 1.960 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 3.625 7.920 5.280 ;
        RECT  4.515 3.705 5.980 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.740 3.700 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.485 -0.400 7.840 1.150 ;
        RECT  4.230 -0.400 4.580 1.035 ;
        RECT  3.500 -0.400 3.840 0.970 ;
        RECT  1.900 -0.400 2.240 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.885 0.620 1.225 ;
        RECT  0.280 0.995 2.460 1.225 ;
        RECT  2.230 1.260 2.645 1.600 ;
        RECT  2.230 0.995 2.460 3.155 ;
        RECT  0.180 2.925 2.460 3.155 ;
        RECT  0.180 2.925 0.520 3.265 ;
        RECT  1.505 2.925 1.845 4.040 ;
        RECT  2.700 0.630 3.160 0.970 ;
        RECT  2.930 0.630 3.160 2.700 ;
        RECT  2.930 2.360 3.825 2.700 ;
        RECT  3.040 2.360 3.305 4.240 ;
        RECT  3.040 3.900 3.380 4.240 ;
        RECT  4.810 0.630 5.355 0.915 ;
        RECT  5.095 0.630 5.355 1.775 ;
        RECT  5.095 1.435 6.515 1.775 ;
        RECT  5.095 0.630 5.325 3.290 ;
        RECT  6.410 2.880 6.750 3.290 ;
        RECT  5.095 2.950 6.750 3.290 ;
        RECT  5.935 0.720 7.060 1.060 ;
        RECT  6.210 3.535 7.200 3.875 ;
        RECT  6.860 3.535 7.200 3.985 ;
        RECT  8.300 0.810 8.640 1.150 ;
        RECT  5.555 2.330 8.640 2.565 ;
        RECT  5.555 2.330 5.840 2.700 ;
        RECT  8.410 0.810 8.640 3.985 ;
        RECT  8.300 3.640 8.640 3.985 ;
        RECT  0.280 0.995 1.30 1.225 ;
        RECT  0.180 2.925 1.70 3.155 ;
        RECT  5.555 2.330 7.10 2.565 ;
    END
END NA6I2X1

MACRO NA6I2X0
    CLASS CORE ;
    FOREIGN NA6I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.250 8.200 2.580 ;
        RECT  7.860 1.955 8.200 2.580 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 3.270 8.695 3.800 ;
        RECT  7.260 3.270 8.695 3.500 ;
        RECT  7.260 2.820 7.550 3.500 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.505 2.675 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.599  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.620 4.105 3.960 ;
        RECT  3.875 1.780 4.105 3.960 ;
        RECT  3.240 1.780 4.105 2.020 ;
        RECT  3.240 1.330 3.655 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 1.990 2.335 ;
        RECT  1.385 2.050 1.765 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.360 1.930 4.915 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.020 4.030 8.360 5.280 ;
        RECT  5.630 3.600 5.970 5.280 ;
        RECT  4.410 3.870 4.750 5.280 ;
        RECT  2.180 3.530 2.520 5.280 ;
        RECT  0.780 3.515 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.170 -0.400 7.510 0.710 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  0.735 1.590 0.965 3.220 ;
        RECT  0.180 2.905 0.965 3.220 ;
        RECT  0.180 2.935 1.710 3.220 ;
        RECT  1.480 2.935 1.710 3.760 ;
        RECT  1.480 3.420 1.820 3.760 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 3.870 ;
        RECT  2.780 2.360 3.645 2.700 ;
        RECT  2.780 2.360 3.045 3.870 ;
        RECT  2.780 3.530 3.335 3.870 ;
        RECT  4.360 0.640 4.700 1.615 ;
        RECT  4.360 1.330 6.380 1.615 ;
        RECT  5.145 1.330 6.380 1.670 ;
        RECT  5.145 1.330 5.375 3.170 ;
        RECT  5.145 2.830 6.570 3.170 ;
        RECT  4.930 2.885 5.270 3.590 ;
        RECT  6.795 1.400 7.510 1.685 ;
        RECT  6.795 1.400 7.030 2.430 ;
        RECT  5.765 2.090 7.030 2.430 ;
        RECT  6.800 1.400 7.030 4.015 ;
        RECT  6.800 3.730 7.285 4.015 ;
        RECT  5.030 0.630 6.825 0.860 ;
        RECT  6.595 0.630 6.825 1.170 ;
        RECT  5.030 0.630 5.370 0.970 ;
        RECT  8.300 0.630 8.660 1.170 ;
        RECT  6.595 0.940 8.660 1.170 ;
        RECT  8.430 0.630 8.660 3.040 ;
        RECT  8.025 2.810 8.660 3.040 ;
        RECT  0.290 1.590 1.30 1.820 ;
        RECT  4.360 1.330 5.20 1.615 ;
        RECT  6.595 0.940 7.80 1.170 ;
    END
END NA6I2X0

MACRO NA6I1X4
    CLASS CORE ;
    FOREIGN NA6I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.145 2.250 8.695 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.881  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.025 3.050 6.825 3.390 ;
        RECT  6.595 1.630 6.825 3.390 ;
        RECT  6.025 1.630 6.825 2.020 ;
        RECT  6.025 1.435 6.370 2.020 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 2.325 2.090 2.710 ;
        RECT  1.435 2.230 1.795 2.710 ;
        END
    END F
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.120 1.600 10.595 2.125 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.220 0.530 3.000 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.865 1.640 1.205 2.540 ;
        RECT  0.735 1.640 1.205 2.035 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.875 7.445 3.240 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.800 3.375 10.155 5.280 ;
        RECT  7.055 4.170 8.515 5.280 ;
        RECT  5.650 3.730 6.015 5.280 ;
        RECT  4.405 3.695 4.745 5.280 ;
        RECT  0.945 4.165 2.405 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.070 -0.400 10.425 1.360 ;
        RECT  6.785 -0.400 7.125 0.710 ;
        RECT  4.995 -0.400 5.335 1.180 ;
        RECT  3.165 -0.400 3.495 0.710 ;
        RECT  1.980 -0.400 2.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.310 0.630 0.650 1.420 ;
        RECT  0.310 1.180 2.310 1.410 ;
        RECT  0.310 1.180 0.655 1.420 ;
        RECT  0.310 0.630 0.640 1.430 ;
        RECT  2.080 1.180 2.310 1.990 ;
        RECT  2.080 1.760 2.875 1.990 ;
        RECT  2.415 1.760 2.875 2.235 ;
        RECT  3.920 2.330 4.505 2.670 ;
        RECT  1.500 2.960 2.875 3.190 ;
        RECT  1.500 2.960 1.845 3.600 ;
        RECT  0.180 3.370 1.845 3.600 ;
        RECT  1.505 2.960 1.845 3.770 ;
        RECT  2.645 1.760 2.875 4.250 ;
        RECT  0.180 3.370 0.535 4.180 ;
        RECT  3.920 2.330 4.175 4.250 ;
        RECT  2.645 4.020 4.175 4.250 ;
        RECT  2.610 1.185 3.495 1.525 ;
        RECT  3.255 1.185 3.495 3.790 ;
        RECT  3.925 1.280 4.270 2.100 ;
        RECT  3.255 1.800 4.270 2.100 ;
        RECT  3.255 1.870 5.595 2.100 ;
        RECT  5.360 1.870 5.595 2.650 ;
        RECT  5.360 2.310 6.365 2.650 ;
        RECT  3.255 1.800 3.620 3.790 ;
        RECT  3.725 0.630 4.735 0.950 ;
        RECT  5.565 0.975 8.835 1.205 ;
        RECT  4.505 0.630 4.735 1.640 ;
        RECT  8.495 0.720 8.835 1.590 ;
        RECT  5.565 0.975 5.795 1.640 ;
        RECT  4.505 1.410 5.795 1.640 ;
        RECT  7.685 0.975 7.915 3.760 ;
        RECT  7.615 3.420 9.275 3.760 ;
        RECT  9.155 1.020 9.605 1.360 ;
        RECT  8.935 2.250 9.385 2.630 ;
        RECT  9.155 1.020 9.385 2.995 ;
        RECT  9.155 2.655 10.155 2.995 ;
        RECT  0.310 1.180 1.60 1.410 ;
        RECT  3.255 1.870 4.60 2.100 ;
        RECT  5.565 0.975 7.90 1.205 ;
    END
END NA6I1X4

MACRO NA6I1X2
    CLASS CORE ;
    FOREIGN NA6I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.530 0.630 2.020 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.675 1.645 8.075 2.165 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.155 1.955 5.510 3.250 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.200 2.195 6.820 2.725 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.685 1.640 4.915 3.360 ;
        RECT  4.475 3.125 4.815 4.045 ;
        RECT  4.535 1.640 4.915 2.020 ;
        RECT  4.190 1.640 4.915 1.870 ;
        RECT  4.190 1.150 4.530 1.870 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.575 1.960 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.360 3.730 7.195 5.280 ;
        RECT  5.235 3.730 5.580 5.280 ;
        RECT  3.715 4.065 4.055 5.280 ;
        RECT  0.885 3.635 2.345 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.865 -0.400 7.210 0.955 ;
        RECT  4.940 -0.400 5.290 1.035 ;
        RECT  3.420 -0.400 3.760 1.220 ;
        RECT  1.900 -0.400 2.240 0.785 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.960 0.620 1.300 ;
        RECT  0.280 1.070 2.460 1.300 ;
        RECT  2.230 1.480 2.660 1.825 ;
        RECT  2.230 1.070 2.460 3.090 ;
        RECT  0.180 2.860 2.460 3.090 ;
        RECT  1.445 2.860 1.785 3.235 ;
        RECT  0.180 2.860 0.520 3.985 ;
        RECT  2.700 0.800 3.160 1.140 ;
        RECT  2.930 0.800 3.160 2.700 ;
        RECT  2.930 2.455 4.455 2.700 ;
        RECT  3.200 2.455 4.455 2.795 ;
        RECT  3.200 2.455 3.540 3.675 ;
        RECT  5.520 0.630 5.985 0.915 ;
        RECT  5.740 0.630 5.985 1.775 ;
        RECT  5.740 1.435 6.985 1.775 ;
        RECT  5.740 0.630 5.970 3.315 ;
        RECT  7.145 2.950 7.485 3.315 ;
        RECT  5.740 2.955 7.485 3.315 ;
        RECT  7.655 0.810 8.010 1.150 ;
        RECT  7.655 0.810 7.930 1.415 ;
        RECT  7.215 1.185 7.930 1.415 ;
        RECT  7.215 1.185 7.445 2.630 ;
        RECT  7.050 2.290 7.445 2.630 ;
        RECT  7.050 2.395 7.945 2.630 ;
        RECT  7.715 2.395 7.945 4.145 ;
        RECT  7.575 3.805 7.945 4.145 ;
        RECT  0.280 1.070 1.80 1.300 ;
        RECT  0.180 2.860 1.20 3.090 ;
    END
END NA6I1X2

MACRO NA6I1X1
    CLASS CORE ;
    FOREIGN NA6I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.505 0.630 2.020 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.105 1.440 7.445 2.095 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.955 4.865 3.240 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.555 2.345 6.125 2.715 ;
        RECT  5.785 2.200 6.125 2.715 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.180 ;
        RECT  3.755 2.930 4.095 3.815 ;
        RECT  3.900 1.640 4.285 2.020 ;
        RECT  3.480 1.640 4.285 1.875 ;
        RECT  3.480 1.480 3.820 1.875 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.495 1.960 2.020 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.840 3.815 6.655 5.280 ;
        RECT  4.515 3.720 4.860 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.740 3.700 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.100 -0.400 6.415 1.020 ;
        RECT  4.230 -0.400 4.580 0.970 ;
        RECT  3.500 -0.400 3.840 0.970 ;
        RECT  1.900 -0.400 2.240 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.885 0.620 1.225 ;
        RECT  0.280 0.995 2.460 1.225 ;
        RECT  2.230 1.260 2.645 1.600 ;
        RECT  2.230 0.995 2.460 3.155 ;
        RECT  0.180 2.925 2.460 3.155 ;
        RECT  0.180 2.925 0.520 3.265 ;
        RECT  1.505 2.925 1.845 4.040 ;
        RECT  2.700 0.630 3.160 0.970 ;
        RECT  2.930 0.630 3.160 4.240 ;
        RECT  2.930 2.360 3.825 2.700 ;
        RECT  2.930 2.360 3.195 4.240 ;
        RECT  2.930 3.900 3.380 4.240 ;
        RECT  4.810 0.630 5.355 0.915 ;
        RECT  5.095 0.630 5.355 1.775 ;
        RECT  5.095 1.435 6.415 1.775 ;
        RECT  5.095 0.630 5.325 3.290 ;
        RECT  6.410 2.890 6.750 3.290 ;
        RECT  5.095 2.950 6.750 3.290 ;
        RECT  6.645 0.770 7.265 1.110 ;
        RECT  6.645 0.770 6.875 2.555 ;
        RECT  6.355 2.215 6.875 2.555 ;
        RECT  6.355 2.325 7.255 2.555 ;
        RECT  7.015 2.325 7.255 4.130 ;
        RECT  7.015 3.790 7.370 4.130 ;
        RECT  0.280 0.995 1.80 1.225 ;
        RECT  0.180 2.925 1.30 3.155 ;
    END
END NA6I1X1

MACRO NA6I1X0
    CLASS CORE ;
    FOREIGN NA6I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.290 1.640 5.575 2.660 ;
        RECT  5.165 1.640 5.575 2.020 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.035 1.475 7.435 2.075 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.505 2.675 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.591  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.600 4.105 3.940 ;
        RECT  3.875 1.785 4.105 3.940 ;
        RECT  3.275 1.785 4.105 2.020 ;
        RECT  3.275 1.330 3.850 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 1.990 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 2.130 4.960 2.660 ;
        RECT  4.520 2.090 4.915 2.660 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.240 3.530 6.580 5.280 ;
        RECT  4.410 3.575 4.750 5.280 ;
        RECT  2.180 3.530 2.520 5.280 ;
        RECT  0.780 3.530 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.240 -0.400 6.580 0.710 ;
        RECT  4.310 -0.400 4.650 1.670 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.180 1.590 2.500 1.820 ;
        RECT  0.735 1.590 0.965 3.220 ;
        RECT  0.180 2.905 0.965 3.220 ;
        RECT  0.180 2.935 1.710 3.220 ;
        RECT  1.480 2.935 1.710 3.760 ;
        RECT  1.480 3.420 1.820 3.760 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 3.870 ;
        RECT  2.780 2.250 3.645 2.590 ;
        RECT  2.780 2.250 3.045 3.870 ;
        RECT  2.780 3.530 3.335 3.870 ;
        RECT  5.670 0.630 6.010 0.915 ;
        RECT  5.780 0.630 6.010 1.470 ;
        RECT  5.805 1.270 6.295 1.620 ;
        RECT  5.805 1.270 6.035 3.220 ;
        RECT  5.805 2.785 6.780 3.070 ;
        RECT  5.010 2.890 6.080 3.220 ;
        RECT  7.040 0.770 7.380 1.170 ;
        RECT  6.525 0.940 7.380 1.170 ;
        RECT  6.265 1.860 6.755 2.205 ;
        RECT  6.525 0.940 6.755 2.555 ;
        RECT  6.525 2.325 7.245 2.555 ;
        RECT  7.015 2.325 7.245 3.870 ;
        RECT  7.015 3.530 7.380 3.870 ;
        RECT  0.180 1.590 1.70 1.820 ;
    END
END NA6I1X0

MACRO NA5X4
    CLASS CORE ;
    FOREIGN NA5X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.250 9.385 2.630 ;
        RECT  9.080 1.900 9.385 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.310 1.640 8.695 2.670 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 3.470 2.150 4.220 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.530 0.525 2.125 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.793  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.400 2.250 7.745 3.920 ;
        RECT  7.245 1.105 7.590 2.630 ;
        RECT  5.960 2.250 7.745 2.630 ;
        RECT  5.960 2.250 6.300 3.920 ;
        RECT  5.960 1.200 6.280 3.920 ;
        RECT  5.805 1.200 6.280 1.580 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  7.965 -0.400 8.305 1.410 ;
        RECT  6.525 -0.400 6.865 1.390 ;
        RECT  5.085 -0.400 5.425 1.445 ;
        RECT  3.605 -0.400 3.945 1.075 ;
        RECT  2.040 -0.400 2.380 1.230 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.560 3.540 9.900 5.280 ;
        RECT  8.120 3.000 8.460 5.280 ;
        RECT  6.680 3.000 7.020 5.280 ;
        RECT  4.680 3.000 5.580 5.280 ;
        RECT  4.680 2.520 5.020 5.280 ;
        RECT  2.380 2.780 2.720 5.280 ;
        RECT  0.900 3.320 1.205 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.420 0.960 1.810 1.300 ;
        RECT  1.580 0.960 1.810 1.745 ;
        RECT  1.790 1.460 2.845 1.820 ;
        RECT  0.180 2.860 2.020 3.090 ;
        RECT  1.790 1.460 2.020 3.145 ;
        RECT  1.620 2.805 2.020 3.145 ;
        RECT  0.180 2.805 0.520 3.700 ;
        RECT  2.845 0.810 3.305 1.150 ;
        RECT  3.075 0.810 3.305 2.165 ;
        RECT  4.365 1.100 4.705 2.170 ;
        RECT  3.075 1.830 5.665 2.165 ;
        RECT  3.530 1.830 5.665 2.170 ;
        RECT  3.530 1.830 3.870 3.840 ;
        RECT  9.560 0.630 9.915 1.545 ;
        RECT  9.145 1.205 9.915 1.545 ;
        RECT  9.615 0.630 9.915 3.230 ;
        RECT  8.840 3.000 9.915 3.230 ;
        RECT  8.840 3.000 9.195 3.920 ;
        RECT  3.075 1.830 4.30 2.165 ;
        RECT  3.530 1.830 4.70 2.170 ;
    END
END NA5X4

MACRO NA5X2
    CLASS CORE ;
    FOREIGN NA5X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.555 1.620 6.865 2.235 ;
        RECT  6.425 1.620 6.865 2.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.770 2.125 6.220 2.470 ;
        RECT  5.770 2.125 6.215 2.670 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.340 3.470 2.060 4.065 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.530 0.525 2.125 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.880 1.225 5.225 3.920 ;
        RECT  4.535 2.250 5.225 2.630 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.600 -0.400 5.940 1.595 ;
        RECT  3.645 -0.400 4.460 1.700 ;
        RECT  2.040 -0.400 2.380 1.230 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 3.080 7.380 5.280 ;
        RECT  5.600 3.050 5.940 5.280 ;
        RECT  4.160 3.000 4.500 5.280 ;
        RECT  2.290 2.780 2.630 5.280 ;
        RECT  0.770 3.595 1.110 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.420 0.960 1.810 1.300 ;
        RECT  1.580 0.960 1.810 1.745 ;
        RECT  1.700 1.460 2.845 1.820 ;
        RECT  1.700 1.460 1.930 3.200 ;
        RECT  0.180 2.860 1.930 3.200 ;
        RECT  2.845 0.810 3.305 1.150 ;
        RECT  3.075 0.810 3.305 2.460 ;
        RECT  3.075 2.125 4.025 2.460 ;
        RECT  3.440 2.125 4.025 2.465 ;
        RECT  3.440 2.125 3.780 4.100 ;
        RECT  7.040 0.630 7.380 1.470 ;
        RECT  7.095 0.630 7.380 2.825 ;
        RECT  6.445 2.595 7.380 2.825 ;
        RECT  6.445 2.595 6.675 3.420 ;
        RECT  6.320 3.080 6.675 3.420 ;
    END
END NA5X2

MACRO NA5X1
    CLASS CORE ;
    FOREIGN NA5X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.430 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.660 3.470 2.395 3.850 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.975 0.525 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.715  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.360 4.380 2.020 ;
        RECT  3.795 3.360 4.135 3.700 ;
        RECT  3.905 1.360 4.135 3.700 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.480 2.240 5.095 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.410 1.640 5.725 2.600 ;
        RECT  5.165 1.640 5.725 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.825 3.600 6.050 5.280 ;
        RECT  2.200 4.080 2.540 5.280 ;
        RECT  0.880 3.595 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.800 -0.400 5.140 0.980 ;
        RECT  3.395 -0.400 3.735 1.105 ;
        RECT  1.790 -0.400 2.130 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.350 2.650 1.690 ;
        RECT  0.290 2.860 1.890 3.090 ;
        RECT  1.660 1.350 1.890 3.200 ;
        RECT  1.440 2.860 1.890 3.200 ;
        RECT  0.290 2.860 0.520 3.940 ;
        RECT  0.180 3.600 0.520 3.940 ;
        RECT  2.595 0.765 3.110 1.105 ;
        RECT  2.880 0.765 3.110 2.490 ;
        RECT  2.880 2.260 3.675 2.490 ;
        RECT  3.190 2.260 3.675 2.600 ;
        RECT  3.190 2.260 3.530 3.120 ;
        RECT  5.780 0.640 6.185 0.980 ;
        RECT  5.150 2.860 6.185 3.090 ;
        RECT  5.955 0.640 6.185 3.090 ;
        RECT  4.365 2.970 5.490 3.200 ;
        RECT  2.950 3.820 3.290 4.160 ;
        RECT  4.365 2.970 4.595 4.160 ;
        RECT  2.950 3.930 4.595 4.160 ;
        RECT  0.180 1.350 1.90 1.690 ;
    END
END NA5X1

MACRO NA5X0
    CLASS CORE ;
    FOREIGN NA5X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.245 0.510 2.875 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.587  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.750 4.135 4.090 ;
        RECT  3.905 1.330 4.135 4.090 ;
        RECT  3.275 1.330 4.135 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.410 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.130 1.900 2.630 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.085 4.940 2.665 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.260 1.540 5.545 2.700 ;
        RECT  5.165 1.540 5.545 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.710 3.730 6.050 5.280 ;
        RECT  4.365 3.080 4.650 5.280 ;
        RECT  2.180 3.730 2.520 5.280 ;
        RECT  0.780 3.730 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.365 -0.400 4.650 1.470 ;
        RECT  3.240 -0.400 4.650 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.870 ;
        RECT  2.160 1.260 2.500 1.870 ;
        RECT  0.290 1.640 2.500 1.870 ;
        RECT  2.215 1.260 2.500 3.365 ;
        RECT  0.180 3.105 2.500 3.365 ;
        RECT  0.180 3.105 1.710 3.420 ;
        RECT  1.480 3.105 1.710 3.960 ;
        RECT  1.480 3.620 1.820 3.960 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 4.070 ;
        RECT  3.360 2.450 3.675 2.790 ;
        RECT  2.780 2.560 3.675 2.790 ;
        RECT  2.780 2.560 3.045 4.070 ;
        RECT  2.780 3.730 3.335 4.070 ;
        RECT  5.720 0.630 6.060 0.950 ;
        RECT  5.750 0.630 6.060 1.435 ;
        RECT  5.775 0.630 6.060 3.420 ;
        RECT  5.110 3.080 6.060 3.420 ;
        RECT  0.290 1.640 1.70 1.870 ;
        RECT  0.180 3.105 1.80 3.365 ;
    END
END NA5X0

MACRO NA5I4X4
    CLASS CORE ;
    FOREIGN NA5I4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.665 2.850 8.065 3.240 ;
        RECT  7.665 2.030 7.895 3.240 ;
        RECT  7.555 2.030 7.895 2.370 ;
        END
    END CN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.240 0.730 2.640 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.940 2.245 9.390 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.260 2.005 8.710 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.881  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.480 3.050 7.270 3.390 ;
        RECT  7.040 1.685 7.270 3.390 ;
        RECT  6.365 1.685 7.270 2.020 ;
        RECT  6.365 1.435 6.805 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.305 2.495 2.730 ;
        RECT  2.005 2.220 2.415 2.730 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.425 3.970 9.770 5.280 ;
        RECT  7.510 4.120 7.855 5.280 ;
        RECT  6.105 3.730 6.470 5.280 ;
        RECT  4.860 3.695 5.200 5.280 ;
        RECT  2.500 4.170 2.840 5.280 ;
        RECT  1.220 3.425 1.560 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  8.885 -0.400 9.710 0.855 ;
        RECT  7.125 -0.400 7.465 0.745 ;
        RECT  5.335 -0.400 5.675 1.180 ;
        RECT  3.530 -0.400 3.860 0.710 ;
        RECT  2.415 -0.400 2.755 0.710 ;
        RECT  0.445 -0.400 0.785 0.900 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.360 0.810 1.855 ;
        RECT  0.445 1.625 1.190 1.855 ;
        RECT  0.960 2.240 1.775 2.580 ;
        RECT  0.960 1.625 1.190 3.105 ;
        RECT  0.460 2.875 1.190 3.105 ;
        RECT  0.460 2.875 0.800 3.215 ;
        RECT  1.220 0.995 1.700 1.335 ;
        RECT  1.470 0.995 1.700 1.990 ;
        RECT  1.470 1.760 3.310 1.990 ;
        RECT  2.780 1.760 3.310 2.235 ;
        RECT  4.270 2.330 4.960 2.670 ;
        RECT  1.940 2.960 3.310 3.190 ;
        RECT  1.940 2.960 2.280 3.770 ;
        RECT  3.080 1.760 3.310 4.250 ;
        RECT  4.270 2.330 4.525 4.250 ;
        RECT  3.080 4.020 4.525 4.250 ;
        RECT  2.975 1.185 3.910 1.525 ;
        RECT  3.680 1.185 3.910 3.790 ;
        RECT  4.290 1.280 4.635 2.100 ;
        RECT  3.680 1.800 4.635 2.100 ;
        RECT  3.680 1.870 6.030 2.100 ;
        RECT  5.795 1.870 6.030 2.650 ;
        RECT  5.795 2.310 6.810 2.650 ;
        RECT  3.680 1.800 4.035 3.790 ;
        RECT  7.910 1.435 8.250 1.775 ;
        RECT  7.910 1.545 9.875 1.775 ;
        RECT  9.380 1.545 9.875 1.995 ;
        RECT  9.645 2.340 10.080 2.680 ;
        RECT  9.645 1.545 9.875 3.425 ;
        RECT  8.930 3.085 9.875 3.425 ;
        RECT  4.090 0.630 5.100 0.915 ;
        RECT  5.905 0.975 8.680 1.205 ;
        RECT  10.125 0.810 10.540 1.315 ;
        RECT  8.480 1.085 10.540 1.315 ;
        RECT  4.870 0.630 5.100 1.640 ;
        RECT  5.905 0.975 6.135 1.640 ;
        RECT  4.870 1.410 6.135 1.640 ;
        RECT  10.310 0.810 10.540 4.165 ;
        RECT  10.190 3.820 10.540 4.165 ;
        RECT  3.680 1.870 5.30 2.100 ;
        RECT  5.905 0.975 7.20 1.205 ;
        RECT  8.480 1.085 9.80 1.315 ;
    END
END NA5I4X4

MACRO NA5I4X2
    CLASS CORE ;
    FOREIGN NA5I4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.885 6.175 3.240 ;
        END
    END CN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.050 2.245 7.500 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.885 6.820 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.315 1.640 5.545 3.395 ;
        RECT  5.015 3.160 5.355 4.080 ;
        RECT  5.150 1.640 5.545 2.020 ;
        RECT  4.800 1.640 5.545 1.870 ;
        RECT  4.800 1.110 5.140 1.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.620 2.405 2.680 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.050 0.540 2.640 ;
        END
    END DN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.535 3.970 7.880 5.280 ;
        RECT  5.775 4.085 6.120 5.280 ;
        RECT  4.290 3.730 4.645 5.280 ;
        RECT  2.475 3.380 2.815 5.280 ;
        RECT  1.030 3.395 1.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.320 -0.400 7.660 0.710 ;
        RECT  5.550 -0.400 5.895 0.970 ;
        RECT  4.010 -0.400 4.350 1.185 ;
        RECT  2.530 -0.400 2.870 0.710 ;
        RECT  0.180 -0.400 0.520 1.025 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.335 1.120 1.680 ;
        RECT  0.780 1.335 1.035 3.100 ;
        RECT  0.780 2.760 1.615 3.100 ;
        RECT  0.425 2.870 1.615 3.100 ;
        RECT  0.425 2.870 0.655 3.700 ;
        RECT  0.315 3.335 0.655 3.700 ;
        RECT  1.300 0.630 1.640 0.980 ;
        RECT  1.400 0.940 2.865 1.170 ;
        RECT  2.635 1.475 3.090 1.830 ;
        RECT  2.635 0.940 2.865 3.140 ;
        RECT  1.865 2.910 2.865 3.140 ;
        RECT  1.865 2.910 2.095 3.740 ;
        RECT  1.750 3.385 2.095 3.740 ;
        RECT  3.290 0.720 3.710 1.060 ;
        RECT  3.480 0.720 3.710 2.585 ;
        RECT  3.620 2.340 5.085 2.680 ;
        RECT  3.620 2.340 3.970 3.365 ;
        RECT  6.200 1.270 6.540 1.630 ;
        RECT  6.200 1.400 7.985 1.630 ;
        RECT  7.600 1.400 7.985 1.785 ;
        RECT  7.755 2.340 8.190 2.680 ;
        RECT  7.755 1.400 7.985 3.395 ;
        RECT  7.195 3.055 7.985 3.395 ;
        RECT  6.125 0.630 7.040 0.915 ;
        RECT  6.810 0.630 7.040 1.170 ;
        RECT  8.140 0.630 8.650 1.170 ;
        RECT  6.810 0.940 8.650 1.170 ;
        RECT  8.420 0.630 8.650 4.135 ;
        RECT  8.300 3.790 8.650 4.135 ;
    END
END NA5I4X2

MACRO NA5I4X1
    CLASS CORE ;
    FOREIGN NA5I4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.560 1.920 4.935 3.240 ;
        END
    END CN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 2.250 2.085 2.670 ;
        END
    END E
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.690 0.505 2.285 ;
        END
    END DN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.790 2.250 6.265 2.780 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.885 5.565 2.200 ;
        RECT  5.165 1.885 5.550 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.772  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.755 2.930 4.330 3.160 ;
        RECT  4.100 1.640 4.330 3.160 ;
        RECT  3.900 1.640 4.330 2.020 ;
        RECT  3.755 2.930 4.095 3.800 ;
        RECT  3.505 1.640 4.330 1.875 ;
        RECT  3.505 1.530 3.850 1.875 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.265 3.970 6.610 5.280 ;
        RECT  4.515 4.085 4.860 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.745 3.790 1.240 5.280 ;
        RECT  0.745 2.975 1.085 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.795 -0.400 6.580 0.710 ;
        RECT  4.265 -0.400 4.595 0.970 ;
        RECT  2.135 -0.400 2.475 0.710 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.170 0.965 1.460 ;
        RECT  0.735 1.680 1.565 2.005 ;
        RECT  0.735 1.170 0.965 2.745 ;
        RECT  0.180 2.515 0.965 2.745 ;
        RECT  0.180 2.515 0.515 4.125 ;
        RECT  1.195 1.110 1.485 1.450 ;
        RECT  1.195 1.205 2.590 1.450 ;
        RECT  2.360 1.855 2.810 2.195 ;
        RECT  2.360 1.205 2.590 3.300 ;
        RECT  1.465 2.960 2.590 3.300 ;
        RECT  2.935 0.630 3.275 0.960 ;
        RECT  3.040 0.630 3.275 4.240 ;
        RECT  3.040 2.360 3.870 2.700 ;
        RECT  3.040 2.360 3.310 4.240 ;
        RECT  3.040 3.900 3.380 4.240 ;
        RECT  4.865 1.310 5.175 1.630 ;
        RECT  4.865 1.325 5.205 1.630 ;
        RECT  4.865 1.400 6.725 1.630 ;
        RECT  6.265 1.400 6.725 1.810 ;
        RECT  6.495 2.340 6.930 2.680 ;
        RECT  6.495 1.400 6.725 3.395 ;
        RECT  5.935 3.055 6.725 3.395 ;
        RECT  4.825 0.630 5.565 0.915 ;
        RECT  5.335 0.630 5.565 1.135 ;
        RECT  7.025 0.630 7.390 1.170 ;
        RECT  5.375 0.940 7.390 1.170 ;
        RECT  7.160 0.630 7.390 4.165 ;
        RECT  7.040 3.820 7.390 4.165 ;
        RECT  5.375 0.940 6.60 1.170 ;
    END
END NA5I4X1

MACRO NA5I4X0
    CLASS CORE ;
    FOREIGN NA5I4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.240 6.225 2.790 ;
        END
    END AN
    PIN DN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.695 2.685 ;
        END
    END DN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.592  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.860 3.620 4.285 3.960 ;
        RECT  4.055 1.640 4.285 3.960 ;
        RECT  3.390 1.640 4.285 2.020 ;
        RECT  3.390 1.330 3.730 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.640 2.145 2.030 ;
        END
    END E
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.860 4.915 3.240 ;
        RECT  4.515 1.865 4.850 3.240 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.860 5.550 2.630 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.925 3.770 7.265 5.280 ;
        RECT  4.560 3.770 4.900 5.280 ;
        RECT  2.330 3.530 2.670 5.280 ;
        RECT  0.930 3.530 1.270 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.760 -0.400 6.575 0.710 ;
        RECT  4.190 -0.400 4.530 0.970 ;
        RECT  3.485 -0.400 3.825 0.970 ;
        RECT  1.885 -0.400 2.230 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.185 1.170 0.525 1.630 ;
        RECT  0.185 1.400 1.155 1.630 ;
        RECT  0.925 2.360 1.620 2.700 ;
        RECT  0.925 1.400 1.155 3.220 ;
        RECT  0.330 2.915 1.155 3.220 ;
        RECT  1.055 0.630 1.395 1.170 ;
        RECT  1.055 0.940 2.385 1.170 ;
        RECT  2.155 1.155 2.700 1.385 ;
        RECT  2.410 1.155 2.700 3.300 ;
        RECT  1.630 3.070 2.700 3.300 ;
        RECT  1.630 3.070 1.970 3.830 ;
        RECT  2.685 0.630 3.160 0.925 ;
        RECT  2.930 0.630 3.160 3.870 ;
        RECT  2.930 2.360 3.825 2.700 ;
        RECT  2.930 2.360 3.195 3.870 ;
        RECT  2.930 3.530 3.485 3.870 ;
        RECT  4.790 1.295 5.105 1.610 ;
        RECT  4.790 1.270 5.075 1.610 ;
        RECT  4.845 1.400 6.800 1.630 ;
        RECT  6.190 1.400 6.800 1.685 ;
        RECT  6.570 1.865 6.985 2.205 ;
        RECT  6.570 1.400 6.800 3.455 ;
        RECT  6.120 3.115 6.800 3.455 ;
        RECT  4.930 0.630 5.530 0.915 ;
        RECT  5.300 0.630 5.530 1.170 ;
        RECT  5.300 0.940 7.445 1.170 ;
        RECT  7.035 0.940 7.445 1.225 ;
        RECT  7.215 0.940 7.445 3.070 ;
        RECT  7.030 2.730 7.445 3.070 ;
        RECT  5.300 0.940 6.40 1.170 ;
    END
END NA5I4X0

MACRO NA5I3X4
    CLASS CORE ;
    FOREIGN NA5I3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 2.245 8.230 3.070 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.995 2.090 7.450 2.635 ;
        END
    END BN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.625 0.515 2.520 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.986  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.850 2.900 6.190 4.180 ;
        RECT  5.780 1.530 6.185 2.030 ;
        RECT  5.780 1.530 6.010 3.390 ;
        RECT  4.490 3.050 6.190 3.390 ;
        RECT  5.265 1.530 6.185 1.780 ;
        RECT  5.265 1.435 5.605 1.780 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.850 6.805 3.240 ;
        RECT  6.425 2.310 6.655 3.240 ;
        RECT  6.295 2.310 6.655 2.650 ;
        END
    END AN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 2.325 1.405 2.710 ;
        RECT  0.745 2.230 1.135 2.710 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.165 3.955 8.510 5.280 ;
        RECT  5.085 3.730 5.450 5.280 ;
        RECT  3.770 3.090 4.110 5.280 ;
        RECT  0.310 4.165 1.770 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.625 -0.400 8.450 0.855 ;
        RECT  6.025 -0.400 6.365 0.745 ;
        RECT  4.235 -0.400 4.575 1.180 ;
        RECT  2.490 -0.400 2.820 0.710 ;
        RECT  1.375 -0.400 1.715 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.010 0.520 1.350 ;
        RECT  0.180 1.120 1.520 1.350 ;
        RECT  1.290 1.120 1.520 1.990 ;
        RECT  1.290 1.760 2.295 1.990 ;
        RECT  1.705 1.760 2.295 2.235 ;
        RECT  3.270 2.330 3.870 2.665 ;
        RECT  0.865 2.960 2.295 3.190 ;
        RECT  0.865 2.960 1.210 3.770 ;
        RECT  2.065 1.760 2.295 4.250 ;
        RECT  3.270 2.330 3.525 4.250 ;
        RECT  2.065 4.020 3.525 4.250 ;
        RECT  1.935 1.185 2.315 1.525 ;
        RECT  1.935 1.280 2.840 1.525 ;
        RECT  2.610 1.280 2.840 3.790 ;
        RECT  3.255 1.280 3.545 2.100 ;
        RECT  2.610 1.830 3.545 2.100 ;
        RECT  2.610 1.870 4.600 2.100 ;
        RECT  4.270 1.870 4.600 2.650 ;
        RECT  4.270 2.310 5.550 2.650 ;
        RECT  2.610 1.830 2.965 3.790 ;
        RECT  6.650 1.435 6.990 1.775 ;
        RECT  6.650 1.545 8.710 1.775 ;
        RECT  8.120 1.545 8.710 1.995 ;
        RECT  8.480 2.200 8.875 2.540 ;
        RECT  8.480 1.545 8.710 3.725 ;
        RECT  6.550 3.470 8.710 3.725 ;
        RECT  6.550 3.470 6.915 3.810 ;
        RECT  3.050 0.630 4.005 0.950 ;
        RECT  4.805 0.975 7.420 1.205 ;
        RECT  8.865 0.810 9.335 1.315 ;
        RECT  7.220 1.085 9.335 1.315 ;
        RECT  3.775 0.630 4.005 1.640 ;
        RECT  4.805 0.975 5.035 1.640 ;
        RECT  3.775 1.410 5.035 1.640 ;
        RECT  9.105 0.810 9.335 4.165 ;
        RECT  8.940 3.240 9.335 4.165 ;
        RECT  6.650 1.545 7.90 1.775 ;
        RECT  6.550 3.470 7.40 3.725 ;
        RECT  4.805 0.975 6.60 1.205 ;
        RECT  7.220 1.085 8.50 1.315 ;
    END
END NA5I3X4

MACRO NA5I3X2
    CLASS CORE ;
    FOREIGN NA5I3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.885 4.915 3.240 ;
        END
    END CN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.790 2.245 6.240 2.785 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.885 5.560 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.395 ;
        RECT  3.755 3.160 4.095 4.080 ;
        RECT  3.540 1.640 4.285 2.020 ;
        RECT  3.540 1.110 3.880 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.640 0.515 2.185 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.235 1.215 2.750 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.275 3.970 6.620 5.280 ;
        RECT  4.515 4.085 4.860 5.280 ;
        RECT  3.030 3.730 3.385 5.280 ;
        RECT  0.175 3.855 1.645 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.060 -0.400 6.400 0.710 ;
        RECT  4.290 -0.400 4.635 0.970 ;
        RECT  2.785 -0.400 3.125 1.355 ;
        RECT  1.270 -0.400 1.610 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.195 1.090 0.535 1.410 ;
        RECT  0.195 1.180 1.675 1.410 ;
        RECT  1.445 1.725 1.890 2.080 ;
        RECT  1.445 1.180 1.675 3.335 ;
        RECT  0.735 3.105 1.675 3.335 ;
        RECT  0.735 3.105 1.080 3.460 ;
        RECT  2.030 0.975 2.450 1.315 ;
        RECT  2.220 0.975 2.450 2.585 ;
        RECT  2.220 2.340 3.825 2.585 ;
        RECT  2.490 2.340 3.825 2.680 ;
        RECT  2.490 2.340 2.840 3.365 ;
        RECT  4.940 1.270 5.280 1.630 ;
        RECT  4.940 1.400 6.725 1.630 ;
        RECT  6.340 1.400 6.725 1.785 ;
        RECT  6.495 2.340 6.930 2.680 ;
        RECT  6.495 1.400 6.725 3.395 ;
        RECT  5.935 3.055 6.725 3.395 ;
        RECT  4.865 0.630 5.780 0.915 ;
        RECT  5.550 0.630 5.780 1.170 ;
        RECT  6.880 0.630 7.390 1.170 ;
        RECT  5.550 0.940 7.390 1.170 ;
        RECT  7.160 0.630 7.390 4.135 ;
        RECT  7.040 3.790 7.390 4.135 ;
    END
END NA5I3X2

MACRO NA5I3X1
    CLASS CORE ;
    FOREIGN NA5I3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.680 0.935 2.020 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.930 1.920 4.295 3.240 ;
        END
    END CN
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.250 1.455 2.670 ;
        END
    END E
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.160 2.250 5.635 2.780 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.211  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.885 4.935 2.200 ;
        RECT  4.535 1.885 4.920 2.630 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.772  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.125 2.930 3.700 3.160 ;
        RECT  3.470 1.635 3.700 3.160 ;
        RECT  2.875 1.635 3.700 2.020 ;
        RECT  3.125 2.930 3.465 3.800 ;
        RECT  2.875 1.530 3.220 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.635 3.970 5.980 5.280 ;
        RECT  3.885 4.085 4.230 5.280 ;
        RECT  1.595 3.900 1.935 5.280 ;
        RECT  0.275 3.700 0.615 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.165 -0.400 5.950 0.710 ;
        RECT  3.635 -0.400 3.965 0.970 ;
        RECT  1.505 -0.400 1.845 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.515 1.110 0.855 1.450 ;
        RECT  0.515 1.205 1.960 1.450 ;
        RECT  1.730 1.855 2.180 2.195 ;
        RECT  1.730 1.205 1.960 3.190 ;
        RECT  0.835 2.960 1.960 3.190 ;
        RECT  0.835 2.960 1.175 3.300 ;
        RECT  2.305 0.630 2.645 0.960 ;
        RECT  2.410 0.630 2.645 4.240 ;
        RECT  2.410 2.360 3.240 2.700 ;
        RECT  2.410 2.360 2.680 4.240 ;
        RECT  2.410 3.900 2.750 4.240 ;
        RECT  4.235 1.305 4.545 1.630 ;
        RECT  4.235 1.325 4.575 1.630 ;
        RECT  4.235 1.400 6.095 1.630 ;
        RECT  5.635 1.400 6.095 1.810 ;
        RECT  5.865 2.340 6.300 2.680 ;
        RECT  5.865 1.400 6.095 3.395 ;
        RECT  5.305 3.055 6.095 3.395 ;
        RECT  4.195 0.630 4.935 0.915 ;
        RECT  4.705 0.630 4.935 1.135 ;
        RECT  6.395 0.630 6.760 1.170 ;
        RECT  4.745 0.940 6.760 1.170 ;
        RECT  6.530 0.630 6.760 4.165 ;
        RECT  6.410 3.820 6.760 4.165 ;
        RECT  4.745 0.940 5.30 1.170 ;
    END
END NA5I3X1

MACRO NA5I3X0
    CLASS CORE ;
    FOREIGN NA5I3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.115 2.205 5.555 2.760 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.215 0.585 3.240 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.593  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.080 3.620 3.475 3.960 ;
        RECT  3.245 1.740 3.475 3.960 ;
        RECT  2.610 1.740 3.475 2.020 ;
        RECT  2.610 1.330 3.025 2.020 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.930 1.640 1.270 2.100 ;
        RECT  0.755 1.640 1.270 2.045 ;
        END
    END E
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.285 3.240 ;
        RECT  3.905 1.890 4.175 3.240 ;
        RECT  3.730 1.890 4.175 2.230 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 1.860 4.885 2.630 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.355 3.440 6.695 5.280 ;
        RECT  3.860 3.770 4.200 5.280 ;
        RECT  1.550 3.530 1.890 5.280 ;
        RECT  0.180 3.770 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.405 -0.400 6.745 0.710 ;
        RECT  5.015 -0.400 5.355 0.710 ;
        RECT  3.410 -0.400 3.750 0.970 ;
        RECT  2.610 -0.400 2.950 0.970 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.870 1.410 ;
        RECT  1.530 1.180 1.870 3.165 ;
        RECT  0.850 2.935 1.870 3.165 ;
        RECT  0.850 2.935 1.190 3.630 ;
        RECT  1.810 0.630 2.380 0.950 ;
        RECT  2.150 0.630 2.380 3.870 ;
        RECT  2.150 2.360 3.015 2.700 ;
        RECT  2.150 2.360 2.415 3.870 ;
        RECT  2.150 3.530 2.705 3.870 ;
        RECT  4.010 1.325 4.370 1.610 ;
        RECT  4.010 1.275 4.350 1.610 ;
        RECT  4.185 1.400 6.125 1.630 ;
        RECT  5.410 1.400 6.125 1.685 ;
        RECT  5.885 1.855 6.200 2.195 ;
        RECT  5.885 1.400 6.125 3.455 ;
        RECT  5.340 3.115 6.125 3.455 ;
        RECT  4.150 0.630 4.785 0.915 ;
        RECT  4.555 0.630 4.785 1.170 ;
        RECT  4.555 0.940 6.745 1.170 ;
        RECT  6.405 0.940 6.745 1.510 ;
        RECT  6.430 0.940 6.745 2.990 ;
        RECT  6.375 2.640 6.745 2.990 ;
        RECT  4.555 0.940 5.40 1.170 ;
    END
END NA5I3X0

MACRO NA5I2X4
    CLASS CORE ;
    FOREIGN NA5I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.835 2.095 8.195 2.460 ;
        RECT  7.685 2.860 8.090 3.245 ;
        RECT  7.835 2.095 8.090 3.245 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.006  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.480 2.970 6.820 4.180 ;
        RECT  6.410 1.530 6.815 2.030 ;
        RECT  6.410 1.530 6.640 3.390 ;
        RECT  5.120 3.050 6.820 3.390 ;
        RECT  5.895 1.530 6.815 1.780 ;
        RECT  5.895 1.435 6.235 1.780 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.700 0.550 3.270 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.920 2.235 7.465 2.680 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 1.625 1.145 2.520 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.325 2.035 2.710 ;
        RECT  1.375 2.230 1.765 2.710 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.165 4.165 8.510 5.280 ;
        RECT  5.715 3.730 6.080 5.280 ;
        RECT  4.400 2.925 4.740 5.280 ;
        RECT  0.940 4.165 2.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.120 -0.400 8.460 0.785 ;
        RECT  6.655 -0.400 6.995 0.745 ;
        RECT  4.865 -0.400 5.205 1.180 ;
        RECT  3.085 -0.400 3.415 0.710 ;
        RECT  1.970 -0.400 2.310 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.340 0.965 0.680 1.395 ;
        RECT  0.340 1.165 2.115 1.395 ;
        RECT  1.885 1.165 2.115 1.990 ;
        RECT  1.885 1.760 2.925 1.990 ;
        RECT  2.335 1.760 2.925 2.235 ;
        RECT  3.900 2.330 4.500 2.665 ;
        RECT  1.495 2.960 2.925 3.190 ;
        RECT  1.495 2.960 1.840 3.770 ;
        RECT  0.180 3.540 1.840 3.770 ;
        RECT  0.180 3.540 0.535 3.900 ;
        RECT  2.695 1.760 2.925 4.250 ;
        RECT  3.900 2.330 4.155 4.250 ;
        RECT  2.695 4.020 4.155 4.250 ;
        RECT  2.530 1.185 2.910 1.525 ;
        RECT  2.530 1.280 3.470 1.525 ;
        RECT  3.240 1.280 3.470 3.790 ;
        RECT  3.850 1.280 4.175 2.100 ;
        RECT  3.240 1.830 4.175 2.100 ;
        RECT  3.240 1.870 5.400 2.100 ;
        RECT  5.165 1.870 5.400 2.650 ;
        RECT  5.165 2.310 6.180 2.650 ;
        RECT  3.240 1.830 3.595 3.790 ;
        RECT  7.280 1.485 7.620 1.825 ;
        RECT  7.280 1.595 8.655 1.825 ;
        RECT  8.425 2.200 8.875 2.540 ;
        RECT  7.180 3.390 7.505 3.730 ;
        RECT  7.180 3.400 7.515 3.730 ;
        RECT  8.425 1.595 8.655 3.730 ;
        RECT  7.180 3.475 8.655 3.730 ;
        RECT  3.645 0.630 4.635 0.950 ;
        RECT  5.435 1.000 8.035 1.205 ;
        RECT  5.435 0.975 7.980 1.205 ;
        RECT  8.875 0.930 9.335 1.360 ;
        RECT  7.815 1.130 9.335 1.360 ;
        RECT  4.405 0.630 4.635 1.640 ;
        RECT  5.435 0.975 5.665 1.640 ;
        RECT  4.405 1.410 5.665 1.640 ;
        RECT  9.105 0.930 9.335 4.045 ;
        RECT  8.930 3.120 9.335 4.045 ;
        RECT  3.240 1.870 4.60 2.100 ;
        RECT  5.435 1.000 7.50 1.205 ;
        RECT  5.435 0.975 6.20 1.205 ;
    END
END NA5I2X4

MACRO NA5I2X2
    CLASS CORE ;
    FOREIGN NA5I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.885 5.545 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.885 6.200 2.630 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 2.200 1.210 2.650 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.685 1.640 4.915 3.395 ;
        RECT  4.385 3.160 4.725 4.080 ;
        RECT  4.520 1.640 4.915 2.020 ;
        RECT  4.170 1.640 4.915 1.870 ;
        RECT  4.170 1.110 4.510 1.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.570 2.285 1.910 2.625 ;
        RECT  1.570 1.620 1.870 2.625 ;
        RECT  1.375 1.620 1.870 2.035 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.425 0.680 1.790 ;
        RECT  0.115 1.425 0.535 2.030 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.315 3.805 6.660 5.280 ;
        RECT  5.145 3.800 5.490 5.280 ;
        RECT  3.660 3.730 4.015 5.280 ;
        RECT  1.890 3.625 2.230 5.280 ;
        RECT  0.180 2.880 0.975 3.225 ;
        RECT  0.180 2.880 0.545 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.600 -0.400 6.940 0.710 ;
        RECT  4.920 -0.400 5.265 0.970 ;
        RECT  3.380 -0.400 3.720 1.185 ;
        RECT  1.900 -0.400 2.240 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.830 0.620 1.170 ;
        RECT  0.280 0.940 2.330 1.170 ;
        RECT  2.100 0.940 2.330 1.830 ;
        RECT  2.230 1.475 2.460 3.115 ;
        RECT  1.240 2.885 2.460 3.115 ;
        RECT  1.240 2.885 1.670 3.225 ;
        RECT  1.240 2.885 1.525 4.145 ;
        RECT  0.895 3.790 1.525 4.145 ;
        RECT  2.690 0.720 3.080 1.060 ;
        RECT  2.850 0.720 3.080 2.585 ;
        RECT  3.075 2.340 4.455 2.680 ;
        RECT  3.075 2.340 3.425 3.365 ;
        RECT  5.570 1.265 5.910 1.630 ;
        RECT  5.570 1.400 6.725 1.630 ;
        RECT  6.495 2.340 6.930 2.680 ;
        RECT  6.495 1.400 6.725 3.395 ;
        RECT  6.135 3.055 6.725 3.395 ;
        RECT  5.495 0.630 6.370 0.915 ;
        RECT  6.140 0.630 6.370 1.170 ;
        RECT  6.140 0.940 7.390 1.170 ;
        RECT  6.975 0.940 7.390 1.700 ;
        RECT  7.160 0.940 7.390 4.150 ;
        RECT  7.040 3.805 7.390 4.150 ;
        RECT  0.280 0.940 1.60 1.170 ;
    END
END NA5I2X2

MACRO NA5I2X1
    CLASS CORE ;
    FOREIGN NA5I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.485 1.875 2.020 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.505 0.630 2.020 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.920 4.915 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.880 5.695 2.630 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.766  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.630 4.285 3.130 ;
        RECT  3.755 2.900 4.095 3.770 ;
        RECT  3.905 1.630 4.285 2.020 ;
        RECT  3.330 1.630 4.285 1.860 ;
        RECT  3.330 1.515 3.640 1.860 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.515 3.800 5.980 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.740 3.700 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.830 -0.400 6.115 0.710 ;
        RECT  4.060 -0.400 4.400 1.400 ;
        RECT  1.800 -0.400 2.140 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.885 0.520 1.225 ;
        RECT  0.180 0.940 2.340 1.225 ;
        RECT  0.180 0.940 1.40 1.225 ;
        RECT  2.110 1.260 2.640 1.600 ;
        RECT  2.110 0.940 2.340 3.210 ;
        RECT  0.180 2.925 2.340 3.210 ;
        RECT  0.180 2.925 1.845 3.265 ;
        RECT  1.505 2.925 1.845 4.040 ;
        RECT  2.600 0.630 3.100 0.950 ;
        RECT  2.870 0.630 3.100 2.670 ;
        RECT  2.870 2.330 3.825 2.670 ;
        RECT  3.130 2.330 3.380 4.240 ;
        RECT  3.040 3.885 3.380 4.240 ;
        RECT  4.860 1.295 5.175 1.630 ;
        RECT  4.860 1.325 5.200 1.630 ;
        RECT  4.860 1.400 6.155 1.630 ;
        RECT  5.925 2.335 6.355 2.675 ;
        RECT  5.925 1.400 6.155 3.240 ;
        RECT  5.650 2.900 6.155 3.240 ;
        RECT  4.795 0.630 5.600 0.915 ;
        RECT  5.370 0.630 5.600 1.170 ;
        RECT  5.370 0.940 6.815 1.170 ;
        RECT  6.385 0.940 6.815 1.465 ;
        RECT  6.585 0.940 6.815 4.185 ;
        RECT  6.410 3.840 6.815 4.185 ;
    END
END NA5I2X1

MACRO NA5I2X0
    CLASS CORE ;
    FOREIGN NA5I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.505 2.675 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.599  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.620 4.135 3.960 ;
        RECT  3.905 1.790 4.135 3.960 ;
        RECT  3.240 1.790 4.135 2.020 ;
        RECT  3.240 1.330 3.655 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 1.990 2.630 ;
        END
    END E
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 2.860 4.915 3.240 ;
        RECT  4.460 2.360 4.870 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.100 2.045 5.495 2.660 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.140 3.440 6.480 5.280 ;
        RECT  4.410 3.530 4.750 5.280 ;
        RECT  2.180 3.530 2.520 5.280 ;
        RECT  0.780 3.530 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.625 -0.400 5.965 0.710 ;
        RECT  4.040 -0.400 4.380 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.290 1.590 2.500 1.820 ;
        RECT  0.735 1.590 0.965 3.220 ;
        RECT  0.180 2.905 0.965 3.220 ;
        RECT  0.180 2.935 1.710 3.220 ;
        RECT  1.480 2.935 1.710 3.760 ;
        RECT  1.480 3.420 1.820 3.760 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 3.870 ;
        RECT  3.360 2.250 3.675 2.590 ;
        RECT  2.780 2.360 3.675 2.590 ;
        RECT  2.780 2.360 3.045 3.870 ;
        RECT  2.780 3.530 3.335 3.870 ;
        RECT  4.740 1.370 5.050 1.670 ;
        RECT  4.740 1.385 5.080 1.670 ;
        RECT  4.740 1.400 5.955 1.670 ;
        RECT  5.725 1.720 6.145 2.060 ;
        RECT  5.725 1.400 5.955 3.245 ;
        RECT  5.350 3.015 5.955 3.245 ;
        RECT  5.350 3.015 5.580 3.870 ;
        RECT  5.240 3.530 5.580 3.870 ;
        RECT  4.660 0.630 5.395 0.915 ;
        RECT  5.165 0.630 5.395 1.170 ;
        RECT  5.165 0.940 6.660 1.170 ;
        RECT  6.320 0.940 6.660 1.510 ;
        RECT  6.375 0.940 6.660 2.980 ;
        RECT  6.185 2.640 6.660 2.980 ;
        RECT  0.290 1.590 1.80 1.820 ;
    END
END NA5I2X0

MACRO NA5I1X4
    CLASS CORE ;
    FOREIGN NA5I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 2.230 2.090 2.710 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.873  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.020 3.050 6.825 3.390 ;
        RECT  6.595 1.630 6.825 3.390 ;
        RECT  6.025 1.630 6.825 2.020 ;
        RECT  6.025 1.435 6.370 2.020 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.840 3.460 9.335 3.955 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.205 2.540 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.220 0.525 3.000 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.205 2.290 7.545 2.660 ;
        RECT  7.055 2.830 7.460 3.240 ;
        RECT  7.205 2.290 7.460 3.240 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.050 4.170 8.510 5.280 ;
        RECT  5.650 3.730 6.015 5.280 ;
        RECT  4.405 3.695 4.745 5.280 ;
        RECT  0.945 4.165 2.405 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.665 -0.400 9.005 0.715 ;
        RECT  6.775 -0.400 7.115 0.710 ;
        RECT  4.995 -0.400 5.335 1.180 ;
        RECT  3.165 -0.400 3.495 0.710 ;
        RECT  1.980 -0.400 2.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.310 0.630 0.650 1.420 ;
        RECT  0.310 1.180 2.310 1.410 ;
        RECT  0.310 1.180 0.655 1.420 ;
        RECT  0.310 0.630 0.640 1.430 ;
        RECT  2.080 1.180 2.310 1.990 ;
        RECT  2.080 1.760 2.875 1.990 ;
        RECT  2.415 1.760 2.875 2.235 ;
        RECT  3.920 2.330 4.505 2.670 ;
        RECT  1.500 2.960 2.875 3.190 ;
        RECT  1.500 2.960 1.845 3.600 ;
        RECT  0.180 3.370 1.845 3.600 ;
        RECT  1.505 2.960 1.845 3.770 ;
        RECT  2.645 1.760 2.875 4.250 ;
        RECT  0.180 3.370 0.535 4.180 ;
        RECT  3.920 2.330 4.175 4.250 ;
        RECT  2.645 4.020 4.175 4.250 ;
        RECT  2.610 1.185 3.495 1.525 ;
        RECT  3.255 1.185 3.495 3.790 ;
        RECT  3.925 1.280 4.270 2.100 ;
        RECT  3.255 1.800 4.270 2.100 ;
        RECT  3.255 1.870 5.595 2.100 ;
        RECT  5.360 1.870 5.595 2.650 ;
        RECT  5.360 2.310 6.365 2.650 ;
        RECT  3.255 1.800 3.620 3.790 ;
        RECT  3.725 0.630 4.735 0.915 ;
        RECT  5.565 0.975 8.305 1.205 ;
        RECT  7.780 0.975 8.305 1.315 ;
        RECT  4.505 0.630 4.735 1.640 ;
        RECT  5.565 0.975 5.795 1.640 ;
        RECT  4.505 1.410 5.795 1.640 ;
        RECT  7.780 0.975 8.010 3.760 ;
        RECT  7.610 3.420 8.010 3.760 ;
        RECT  8.240 1.865 9.005 2.210 ;
        RECT  8.660 1.170 9.005 3.220 ;
        RECT  8.655 1.865 9.005 3.220 ;
        RECT  8.655 2.880 9.275 3.220 ;
        RECT  0.310 1.180 1.80 1.410 ;
        RECT  3.255 1.870 4.70 2.100 ;
        RECT  5.565 0.975 7.00 1.205 ;
    END
END NA5I1X4

MACRO NA5I1X2
    CLASS CORE ;
    FOREIGN NA5I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.360 1.550 1.890 2.020 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.435 2.630 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.045 2.305 7.445 2.820 ;
        RECT  7.065 2.245 7.445 2.820 ;
        RECT  7.060 2.255 7.445 2.820 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.530 0.630 2.020 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.163  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.155 2.090 5.510 3.250 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.685 1.640 4.915 3.360 ;
        RECT  4.455 3.125 4.795 4.045 ;
        RECT  4.535 1.640 4.915 2.020 ;
        RECT  4.095 1.640 4.915 1.870 ;
        RECT  4.095 1.150 4.435 1.870 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.200 3.050 7.445 5.280 ;
        RECT  6.755 3.050 7.445 3.390 ;
        RECT  5.175 3.610 5.520 5.280 ;
        RECT  3.695 4.065 4.035 5.280 ;
        RECT  0.885 3.635 2.345 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.235 -0.400 6.580 0.955 ;
        RECT  4.845 -0.400 5.195 1.035 ;
        RECT  3.325 -0.400 3.665 1.220 ;
        RECT  1.805 -0.400 2.145 0.785 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.185 0.960 0.525 1.300 ;
        RECT  0.185 1.070 2.365 1.300 ;
        RECT  2.135 1.070 2.365 3.090 ;
        RECT  2.135 1.480 2.565 1.825 ;
        RECT  2.135 1.480 2.460 3.090 ;
        RECT  0.180 2.860 2.460 3.090 ;
        RECT  1.445 2.860 1.785 3.235 ;
        RECT  0.180 2.860 0.520 3.985 ;
        RECT  2.605 0.800 3.065 1.140 ;
        RECT  2.835 0.800 3.065 2.755 ;
        RECT  2.835 2.510 4.455 2.755 ;
        RECT  3.195 2.510 4.455 2.850 ;
        RECT  3.195 2.510 3.535 3.675 ;
        RECT  5.425 0.630 5.985 0.915 ;
        RECT  5.740 0.630 5.985 1.775 ;
        RECT  5.740 1.435 6.400 1.775 ;
        RECT  5.740 0.630 5.970 3.125 ;
        RECT  5.740 2.765 6.065 3.125 ;
        RECT  7.040 0.810 7.380 1.435 ;
        RECT  6.630 1.205 7.380 1.435 ;
        RECT  6.630 1.205 6.860 2.140 ;
        RECT  6.200 2.005 6.825 2.235 ;
        RECT  6.200 2.005 6.545 2.365 ;
        RECT  6.295 2.005 6.525 4.250 ;
        RECT  6.295 3.930 6.970 4.250 ;
        RECT  0.185 1.070 1.60 1.300 ;
        RECT  0.180 2.860 1.50 3.090 ;
    END
END NA5I1X2

MACRO NA5I1X1
    CLASS CORE ;
    FOREIGN NA5I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.495 1.960 2.020 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.530 2.630 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.370 2.300 6.815 2.755 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.505 0.630 2.020 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.955 4.865 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.160 ;
        RECT  3.755 2.930 4.095 3.815 ;
        RECT  3.480 1.640 4.285 2.020 ;
        RECT  3.480 1.480 3.820 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.515 3.715 5.985 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.740 3.700 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.585 -0.400 5.930 0.970 ;
        RECT  4.230 -0.400 4.580 1.055 ;
        RECT  3.500 -0.400 3.840 0.970 ;
        RECT  1.900 -0.400 2.240 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 0.885 0.620 1.225 ;
        RECT  0.280 0.940 2.460 1.225 ;
        RECT  2.230 1.260 2.645 1.600 ;
        RECT  2.230 0.940 2.460 3.210 ;
        RECT  0.180 2.925 2.460 3.210 ;
        RECT  0.180 2.925 1.845 3.265 ;
        RECT  1.505 2.925 1.845 4.040 ;
        RECT  2.700 0.630 3.160 0.970 ;
        RECT  2.930 0.630 3.160 4.240 ;
        RECT  2.930 2.360 3.825 2.700 ;
        RECT  2.930 2.360 3.195 4.240 ;
        RECT  2.930 3.900 3.380 4.240 ;
        RECT  4.810 0.630 5.355 0.915 ;
        RECT  5.095 0.630 5.355 1.625 ;
        RECT  5.095 1.330 5.925 1.625 ;
        RECT  5.095 0.630 5.325 3.290 ;
        RECT  5.095 2.950 5.415 3.290 ;
        RECT  6.410 0.720 6.750 1.060 ;
        RECT  6.015 1.840 6.640 2.070 ;
        RECT  6.410 0.720 6.640 2.070 ;
        RECT  5.560 2.010 6.140 2.350 ;
        RECT  5.910 1.855 6.140 3.270 ;
        RECT  5.910 2.985 6.740 3.270 ;
        RECT  0.280 0.940 1.60 1.225 ;
        RECT  0.180 2.925 1.60 3.210 ;
    END
END NA5I1X1

MACRO NA5I1X0
    CLASS CORE ;
    FOREIGN NA5I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.075 0.505 2.675 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.599  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 3.620 4.135 3.960 ;
        RECT  3.905 1.790 4.135 3.960 ;
        RECT  3.240 1.790 4.135 2.020 ;
        RECT  3.240 1.330 3.655 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.050 2.000 2.630 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 2.050 4.870 2.700 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.180 2.280 6.805 2.675 ;
        RECT  6.425 2.250 6.805 2.675 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.410 3.580 5.950 5.280 ;
        RECT  2.180 3.530 2.520 5.280 ;
        RECT  0.780 3.530 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.870 -0.400 6.210 0.710 ;
        RECT  4.040 -0.400 4.380 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.820 ;
        RECT  2.160 1.260 2.500 1.820 ;
        RECT  0.180 1.590 2.500 1.820 ;
        RECT  0.735 1.590 0.965 3.220 ;
        RECT  0.180 2.905 0.965 3.220 ;
        RECT  0.180 2.935 1.710 3.220 ;
        RECT  1.480 2.935 1.710 3.760 ;
        RECT  1.480 3.420 1.820 3.760 ;
        RECT  2.440 0.630 3.010 0.970 ;
        RECT  2.780 0.630 3.010 3.870 ;
        RECT  3.360 2.250 3.675 2.590 ;
        RECT  2.780 2.360 3.675 2.590 ;
        RECT  2.780 2.360 3.045 3.870 ;
        RECT  2.780 3.530 3.335 3.870 ;
        RECT  4.660 0.630 5.330 0.915 ;
        RECT  5.100 1.170 5.510 1.510 ;
        RECT  5.100 0.630 5.330 3.220 ;
        RECT  5.065 2.880 5.330 3.220 ;
        RECT  5.010 2.885 5.335 3.220 ;
        RECT  5.870 1.170 6.210 2.050 ;
        RECT  5.560 1.820 6.210 2.050 ;
        RECT  5.560 1.820 5.850 2.270 ;
        RECT  5.565 1.820 5.850 3.165 ;
        RECT  5.565 2.905 6.750 3.165 ;
        RECT  6.410 2.905 6.750 3.220 ;
        RECT  0.180 1.590 1.30 1.820 ;
    END
END NA5I1X0

MACRO NA4X4
    CLASS CORE ;
    FOREIGN NA4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.415 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.650 2.245 8.145 2.630 ;
        RECT  7.650 2.125 8.110 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.575 0.525 2.175 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.565 1.700 8.875 2.270 ;
        RECT  8.315 1.620 8.745 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.793  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.720 1.640 7.435 2.020 ;
        RECT  6.725 1.175 7.070 3.745 ;
        RECT  5.275 2.025 7.070 2.255 ;
        RECT  6.720 1.175 7.070 2.255 ;
        RECT  5.275 1.200 5.625 3.745 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.930 2.960 9.270 5.280 ;
        RECT  7.450 2.860 7.790 5.280 ;
        RECT  6.005 2.825 6.345 5.280 ;
        RECT  3.920 2.730 4.865 5.280 ;
        RECT  4.525 2.680 4.865 5.280 ;
        RECT  1.620 3.540 1.960 5.280 ;
        RECT  0.180 3.075 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.445 -0.400 7.785 1.410 ;
        RECT  6.005 -0.400 6.345 1.540 ;
        RECT  4.565 -0.400 4.905 1.410 ;
        RECT  2.770 -0.400 3.110 1.115 ;
        RECT  1.330 -0.400 1.670 1.060 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.800 0.520 1.220 ;
        RECT  0.180 0.935 1.030 1.220 ;
        RECT  0.800 0.935 1.030 1.575 ;
        RECT  0.800 1.290 1.845 1.575 ;
        RECT  1.615 1.540 2.070 1.660 ;
        RECT  1.645 1.540 2.070 1.880 ;
        RECT  3.345 2.160 4.020 2.500 ;
        RECT  1.645 1.540 1.875 3.310 ;
        RECT  0.900 3.080 2.540 3.310 ;
        RECT  0.900 3.080 1.240 4.000 ;
        RECT  2.310 3.080 2.540 4.250 ;
        RECT  3.345 2.160 3.575 4.250 ;
        RECT  2.310 4.020 3.575 4.250 ;
        RECT  2.050 0.815 2.540 1.155 ;
        RECT  2.310 0.815 2.540 1.595 ;
        RECT  2.310 1.365 4.335 1.595 ;
        RECT  3.530 1.310 4.335 1.650 ;
        RECT  2.770 1.365 4.335 1.650 ;
        RECT  4.105 1.700 4.495 1.935 ;
        RECT  4.105 1.310 4.335 1.935 ;
        RECT  4.250 1.900 5.045 2.240 ;
        RECT  2.770 1.365 3.115 3.790 ;
        RECT  8.930 0.630 9.335 1.470 ;
        RECT  9.105 0.630 9.335 2.730 ;
        RECT  8.470 2.500 9.335 2.730 ;
        RECT  8.470 2.500 8.700 3.245 ;
        RECT  8.210 2.905 8.700 3.245 ;
        RECT  2.310 1.365 3.20 1.595 ;
    END
END NA4X4

MACRO NA4X2
    CLASS CORE ;
    FOREIGN NA4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.415 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.140 2.125 5.590 2.470 ;
        RECT  5.140 2.125 5.585 2.670 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.235 0.520 2.845 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.925 1.620 6.235 2.235 ;
        RECT  5.795 1.620 6.235 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.320 1.640 4.915 2.020 ;
        RECT  4.190 3.000 4.550 3.920 ;
        RECT  4.320 1.175 4.550 3.920 ;
        RECT  4.200 1.175 4.550 1.515 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.080 6.750 5.280 ;
        RECT  4.930 3.000 5.270 5.280 ;
        RECT  3.485 3.000 3.825 5.280 ;
        RECT  1.500 3.820 1.840 5.280 ;
        RECT  0.180 3.075 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.000 -0.400 5.340 1.410 ;
        RECT  2.815 -0.400 3.825 1.650 ;
        RECT  1.210 -0.400 1.550 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.350 0.520 1.825 ;
        RECT  0.180 1.540 2.070 1.825 ;
        RECT  1.645 1.540 2.070 1.880 ;
        RECT  1.645 1.540 1.875 3.380 ;
        RECT  0.900 3.040 1.875 3.380 ;
        RECT  2.015 0.815 2.585 1.155 ;
        RECT  2.355 0.815 2.585 2.235 ;
        RECT  2.355 1.900 3.305 2.235 ;
        RECT  2.690 1.900 3.305 2.240 ;
        RECT  2.690 1.900 3.030 4.000 ;
        RECT  6.410 0.630 6.750 1.470 ;
        RECT  6.465 0.630 6.750 2.825 ;
        RECT  5.815 2.595 6.750 2.825 ;
        RECT  5.815 2.595 6.045 3.420 ;
        RECT  5.690 3.080 6.045 3.420 ;
    END
END NA4X2

MACRO NA4X1
    CLASS CORE ;
    FOREIGN NA4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.130 0.800 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.960 3.470 1.765 3.850 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.715  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.410 1.360 3.750 2.020 ;
        RECT  3.165 3.360 3.505 3.700 ;
        RECT  3.275 1.640 3.505 3.700 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.850 2.240 4.465 2.635 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.780 2.260 5.095 2.600 ;
        RECT  4.780 1.640 5.010 2.600 ;
        RECT  4.535 1.640 5.010 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.195 3.600 5.420 5.280 ;
        RECT  1.500 4.080 1.840 5.280 ;
        RECT  0.180 3.595 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.170 -0.400 4.510 0.980 ;
        RECT  2.775 -0.400 3.115 1.095 ;
        RECT  1.170 -0.400 1.510 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.350 2.030 1.690 ;
        RECT  1.030 1.350 1.260 3.200 ;
        RECT  0.740 2.860 1.260 3.200 ;
        RECT  1.975 0.755 2.490 1.095 ;
        RECT  2.260 0.755 2.490 2.490 ;
        RECT  2.490 2.260 3.045 2.600 ;
        RECT  2.490 2.260 2.830 3.120 ;
        RECT  5.150 0.640 5.555 0.980 ;
        RECT  4.520 2.860 5.555 3.090 ;
        RECT  5.325 0.640 5.555 3.090 ;
        RECT  3.735 2.970 4.860 3.200 ;
        RECT  2.250 3.820 2.590 4.160 ;
        RECT  3.735 2.970 3.965 4.160 ;
        RECT  2.250 3.930 3.965 4.160 ;
    END
END NA4X1

MACRO NA4X0
    CLASS CORE ;
    FOREIGN NA4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.505 2.900 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.587  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.655 2.020 ;
        RECT  3.110 3.930 3.505 4.250 ;
        RECT  3.275 1.330 3.505 4.250 ;
        RECT  2.905 1.330 3.505 1.670 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.415 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 2.130 4.330 2.660 ;
        RECT  3.890 2.090 4.285 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.690 1.640 4.975 3.100 ;
        RECT  4.535 1.640 4.975 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 3.820 5.490 5.280 ;
        RECT  3.740 3.280 4.080 5.280 ;
        RECT  1.580 3.930 1.920 5.280 ;
        RECT  0.180 3.275 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.740 -0.400 4.080 1.380 ;
        RECT  2.815 -0.400 4.080 0.970 ;
        RECT  1.210 -0.400 1.550 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.520 1.510 ;
        RECT  0.180 1.225 2.015 1.510 ;
        RECT  1.645 1.225 2.015 1.565 ;
        RECT  1.645 1.225 1.875 3.565 ;
        RECT  0.880 3.335 1.875 3.565 ;
        RECT  0.880 3.335 1.110 4.230 ;
        RECT  0.880 3.890 1.220 4.230 ;
        RECT  2.015 0.630 2.475 0.970 ;
        RECT  2.245 2.670 3.045 3.030 ;
        RECT  2.245 0.630 2.475 4.250 ;
        RECT  2.245 3.930 2.735 4.250 ;
        RECT  5.150 0.630 5.490 1.470 ;
        RECT  5.205 0.630 5.490 3.565 ;
        RECT  4.550 3.335 5.490 3.565 ;
        RECT  4.550 3.335 4.780 4.250 ;
        RECT  4.440 3.930 4.780 4.250 ;
    END
END NA4X0

MACRO NA4I3X4
    CLASS CORE ;
    FOREIGN NA4I3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.240 0.730 2.640 ;
        END
    END CN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 2.305 2.495 2.730 ;
        RECT  2.005 2.220 2.415 2.730 ;
        END
    END D
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.295 2.195 8.710 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.545 2.230 8.065 2.700 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.928  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.580 3.050 7.270 3.390 ;
        RECT  7.040 1.685 7.270 3.390 ;
        RECT  6.365 1.685 7.270 2.020 ;
        RECT  6.365 1.435 6.805 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.795 3.970 9.140 5.280 ;
        RECT  6.210 3.730 6.550 5.280 ;
        RECT  4.860 3.070 5.200 5.280 ;
        RECT  2.500 4.170 2.840 5.280 ;
        RECT  1.220 3.425 1.560 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.780 -0.400 9.120 1.010 ;
        RECT  7.125 -0.400 7.465 0.745 ;
        RECT  5.335 -0.400 5.675 1.180 ;
        RECT  2.415 -0.400 3.860 0.710 ;
        RECT  0.445 -0.400 0.785 0.900 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.360 0.810 1.855 ;
        RECT  0.445 1.625 1.190 1.855 ;
        RECT  0.960 2.240 1.775 2.580 ;
        RECT  0.960 1.625 1.190 3.105 ;
        RECT  0.460 2.875 1.190 3.105 ;
        RECT  0.460 2.875 0.800 3.215 ;
        RECT  1.220 0.995 1.700 1.335 ;
        RECT  1.470 0.995 1.700 1.990 ;
        RECT  1.470 1.760 3.310 1.990 ;
        RECT  2.780 1.760 3.310 2.235 ;
        RECT  4.270 2.330 4.960 2.665 ;
        RECT  1.940 2.960 3.310 3.190 ;
        RECT  1.940 2.960 2.280 3.770 ;
        RECT  3.080 1.760 3.310 4.250 ;
        RECT  4.270 2.330 4.525 4.250 ;
        RECT  3.080 4.020 4.525 4.250 ;
        RECT  2.975 1.185 3.910 1.525 ;
        RECT  3.680 1.185 3.910 3.790 ;
        RECT  4.290 1.280 4.635 2.100 ;
        RECT  3.680 1.800 4.635 2.100 ;
        RECT  3.680 1.870 5.595 2.100 ;
        RECT  5.360 1.870 5.595 2.650 ;
        RECT  5.360 2.310 6.810 2.650 ;
        RECT  3.680 1.800 4.035 3.790 ;
        RECT  7.790 1.600 8.130 1.940 ;
        RECT  7.790 1.700 9.245 1.940 ;
        RECT  9.015 2.340 9.405 2.680 ;
        RECT  7.610 3.330 7.950 3.700 ;
        RECT  9.015 1.700 9.245 3.700 ;
        RECT  7.610 3.470 9.245 3.700 ;
        RECT  4.090 0.630 5.100 0.915 ;
        RECT  5.905 0.975 8.550 1.205 ;
        RECT  8.320 0.975 8.550 1.470 ;
        RECT  4.870 0.630 5.100 1.640 ;
        RECT  9.540 1.130 9.910 1.470 ;
        RECT  8.320 1.240 9.910 1.470 ;
        RECT  5.905 0.975 6.135 1.640 ;
        RECT  4.870 1.410 6.135 1.640 ;
        RECT  9.680 1.130 9.910 4.090 ;
        RECT  9.560 3.745 9.910 4.090 ;
        RECT  5.905 0.975 7.40 1.205 ;
    END
END NA4I3X4

MACRO NA4I3X2
    CLASS CORE ;
    FOREIGN NA4I3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.050 0.540 2.640 ;
        END
    END CN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 1.925 6.175 3.240 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.940 3.160 5.545 3.395 ;
        RECT  5.315 1.640 5.545 3.395 ;
        RECT  5.150 1.640 5.545 2.020 ;
        RECT  4.940 3.160 5.280 4.080 ;
        RECT  4.800 1.640 5.545 1.870 ;
        RECT  4.800 1.110 5.140 1.870 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.415 2.045 6.830 2.640 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.620 2.405 2.035 ;
        RECT  1.995 1.620 2.335 2.680 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  5.700 3.825 7.250 5.280 ;
        RECT  4.215 3.730 4.570 5.280 ;
        RECT  2.475 3.380 2.815 5.280 ;
        RECT  1.030 3.395 1.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.230 -0.400 7.570 0.710 ;
        RECT  5.550 -0.400 5.895 0.970 ;
        RECT  4.010 -0.400 4.350 1.185 ;
        RECT  2.530 -0.400 2.870 0.710 ;
        RECT  0.180 -0.400 0.520 1.025 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 1.335 1.120 3.100 ;
        RECT  0.780 2.760 1.615 3.100 ;
        RECT  0.315 2.870 1.615 3.100 ;
        RECT  0.315 2.870 0.655 3.700 ;
        RECT  1.300 0.630 1.640 0.980 ;
        RECT  1.400 0.940 2.865 1.170 ;
        RECT  2.635 1.475 3.090 1.830 ;
        RECT  2.635 0.940 2.865 3.140 ;
        RECT  1.865 2.910 2.865 3.140 ;
        RECT  1.865 2.910 2.095 3.740 ;
        RECT  1.750 3.385 2.095 3.740 ;
        RECT  3.290 0.720 3.710 1.060 ;
        RECT  3.480 0.720 3.710 2.585 ;
        RECT  3.620 2.340 5.085 2.680 ;
        RECT  3.620 2.340 3.970 3.365 ;
        RECT  6.200 1.270 6.540 1.630 ;
        RECT  6.200 1.400 7.320 1.630 ;
        RECT  7.090 2.340 7.495 2.680 ;
        RECT  7.090 1.400 7.320 3.270 ;
        RECT  6.690 2.930 7.320 3.270 ;
        RECT  6.125 0.630 7.000 0.915 ;
        RECT  6.770 0.630 7.000 1.170 ;
        RECT  6.770 0.940 7.895 1.170 ;
        RECT  7.665 0.940 7.895 1.700 ;
        RECT  7.790 1.345 8.020 4.135 ;
        RECT  7.670 3.790 8.020 4.135 ;
    END
END NA4I3X2

MACRO NA4I3X1
    CLASS CORE ;
    FOREIGN NA4I3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.690 0.505 2.285 ;
        END
    END CN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 2.250 2.085 2.670 ;
        END
    END D
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.560 1.920 4.925 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.885 5.605 2.630 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.772  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.755 2.930 4.330 3.160 ;
        RECT  4.100 1.640 4.330 3.160 ;
        RECT  3.505 1.640 4.330 2.020 ;
        RECT  3.755 2.930 4.095 3.800 ;
        RECT  3.505 1.530 3.845 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.685 3.800 6.030 5.280 ;
        RECT  4.515 3.900 4.860 5.280 ;
        RECT  2.225 3.900 2.565 5.280 ;
        RECT  0.745 3.790 1.240 5.280 ;
        RECT  0.745 2.975 1.085 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.795 -0.400 6.080 0.710 ;
        RECT  4.265 -0.400 4.595 0.970 ;
        RECT  2.135 -0.400 2.475 0.710 ;
        RECT  0.445 -0.400 0.785 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.170 0.965 1.460 ;
        RECT  0.735 1.680 1.565 2.005 ;
        RECT  0.735 1.170 0.965 2.745 ;
        RECT  0.180 2.515 0.965 2.745 ;
        RECT  0.180 2.515 0.515 4.125 ;
        RECT  1.195 1.110 1.485 1.450 ;
        RECT  1.195 1.205 2.590 1.450 ;
        RECT  2.360 1.855 2.810 2.195 ;
        RECT  2.360 1.205 2.590 3.190 ;
        RECT  1.465 2.960 2.590 3.190 ;
        RECT  1.465 2.960 1.805 3.300 ;
        RECT  2.935 0.630 3.275 0.960 ;
        RECT  3.040 0.630 3.275 4.240 ;
        RECT  3.040 2.360 3.870 2.700 ;
        RECT  3.040 2.360 3.310 4.240 ;
        RECT  3.040 3.900 3.380 4.240 ;
        RECT  4.865 1.305 5.175 1.630 ;
        RECT  4.865 1.325 5.205 1.630 ;
        RECT  4.865 1.400 6.095 1.630 ;
        RECT  5.865 2.205 6.280 2.545 ;
        RECT  5.865 1.400 6.095 3.220 ;
        RECT  5.675 2.880 6.095 3.220 ;
        RECT  4.825 0.630 5.565 0.915 ;
        RECT  5.335 0.630 5.565 1.135 ;
        RECT  5.375 0.940 6.760 1.170 ;
        RECT  6.410 0.940 6.760 1.360 ;
        RECT  6.530 0.940 6.760 4.150 ;
        RECT  6.410 3.805 6.760 4.150 ;
    END
END NA4I3X1

MACRO NA4I3X0
    CLASS CORE ;
    FOREIGN NA4I3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.745 2.630 ;
        RECT  0.440 2.060 0.745 2.630 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.285 2.020 ;
        RECT  3.740 3.620 4.135 3.960 ;
        RECT  3.905 1.330 4.135 3.960 ;
        RECT  3.445 1.330 4.135 1.670 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 1.755 2.115 2.095 ;
        RECT  1.435 1.640 1.765 2.095 ;
        END
    END D
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.500 2.105 4.935 2.650 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.360 5.605 3.240 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.440 6.750 5.280 ;
        RECT  4.370 2.880 4.710 5.280 ;
        RECT  2.210 3.530 2.550 5.280 ;
        RECT  0.810 3.525 1.150 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.730 -0.400 6.070 0.710 ;
        RECT  4.245 -0.400 4.590 0.970 ;
        RECT  3.515 -0.400 3.855 0.970 ;
        RECT  1.910 -0.400 2.250 0.710 ;
        RECT  0.210 -0.400 0.550 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.210 1.170 0.550 1.630 ;
        RECT  0.210 1.400 1.205 1.630 ;
        RECT  0.975 2.360 1.520 2.700 ;
        RECT  0.975 1.400 1.205 3.220 ;
        RECT  0.180 2.880 1.205 3.220 ;
        RECT  1.080 0.630 1.420 1.170 ;
        RECT  1.080 0.940 2.415 1.170 ;
        RECT  2.185 1.145 2.715 1.430 ;
        RECT  2.345 1.145 2.715 1.490 ;
        RECT  2.345 1.145 2.575 3.165 ;
        RECT  1.510 2.935 2.575 3.165 ;
        RECT  1.510 2.935 1.740 3.830 ;
        RECT  1.510 3.490 1.850 3.830 ;
        RECT  2.715 0.630 3.175 0.915 ;
        RECT  2.945 0.630 3.175 2.700 ;
        RECT  2.875 2.360 3.675 2.700 ;
        RECT  2.875 2.360 3.105 3.870 ;
        RECT  2.875 3.530 3.365 3.870 ;
        RECT  4.805 1.370 5.155 1.670 ;
        RECT  4.805 1.385 5.185 1.670 ;
        RECT  4.805 1.400 6.065 1.670 ;
        RECT  5.835 1.785 6.330 2.100 ;
        RECT  5.835 1.400 6.065 3.870 ;
        RECT  5.400 3.530 6.065 3.870 ;
        RECT  4.820 0.630 5.500 0.915 ;
        RECT  5.270 0.630 5.500 1.170 ;
        RECT  5.270 0.940 6.675 1.170 ;
        RECT  6.320 0.940 6.675 1.485 ;
        RECT  6.585 1.240 6.815 2.980 ;
        RECT  6.295 2.640 6.815 2.980 ;
    END
END NA4I3X0

MACRO NA4I2X4
    CLASS CORE ;
    FOREIGN NA4I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 2.230 1.275 2.710 ;
        END
    END D
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.035 2.195 7.450 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.325 2.215 6.805 2.720 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.973  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 1.630 6.185 2.030 ;
        RECT  4.380 3.050 6.010 3.390 ;
        RECT  5.780 1.630 6.010 3.390 ;
        RECT  5.290 1.630 6.185 1.880 ;
        RECT  5.290 1.435 5.635 1.880 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.200 0.515 2.810 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.535 3.970 7.880 5.280 ;
        RECT  5.010 3.730 5.350 5.280 ;
        RECT  3.660 2.930 4.000 5.280 ;
        RECT  0.180 4.165 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.520 -0.400 7.860 0.970 ;
        RECT  6.050 -0.400 6.390 0.745 ;
        RECT  4.260 -0.400 4.600 1.180 ;
        RECT  1.370 -0.400 2.815 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 1.550 1.510 ;
        RECT  1.320 1.170 1.550 1.990 ;
        RECT  1.320 1.760 2.105 1.990 ;
        RECT  1.685 1.760 2.105 2.235 ;
        RECT  3.060 2.330 3.785 2.665 ;
        RECT  0.740 2.960 2.105 3.190 ;
        RECT  0.740 2.960 1.080 3.770 ;
        RECT  1.875 1.760 2.105 4.250 ;
        RECT  3.060 2.330 3.315 4.250 ;
        RECT  1.875 4.020 3.315 4.250 ;
        RECT  1.930 1.185 2.710 1.525 ;
        RECT  2.480 1.185 2.710 3.790 ;
        RECT  3.245 1.280 3.570 2.100 ;
        RECT  2.480 1.800 3.570 2.100 ;
        RECT  2.480 1.870 4.395 2.100 ;
        RECT  4.160 1.870 4.395 2.650 ;
        RECT  4.160 2.310 5.550 2.650 ;
        RECT  2.480 1.800 2.830 3.790 ;
        RECT  6.650 1.600 6.990 1.940 ;
        RECT  6.650 1.700 7.985 1.940 ;
        RECT  7.755 2.340 8.145 2.680 ;
        RECT  6.350 3.330 6.690 3.700 ;
        RECT  7.755 1.700 7.985 3.700 ;
        RECT  6.350 3.470 7.985 3.700 ;
        RECT  3.045 0.630 4.030 0.915 ;
        RECT  4.830 0.975 7.290 1.205 ;
        RECT  7.060 1.200 8.650 1.380 ;
        RECT  3.800 0.630 4.030 1.640 ;
        RECT  7.145 1.200 8.650 1.430 ;
        RECT  8.280 1.130 8.650 1.470 ;
        RECT  4.830 0.975 5.060 1.640 ;
        RECT  3.800 1.410 5.060 1.640 ;
        RECT  8.420 1.130 8.650 4.090 ;
        RECT  8.300 3.165 8.650 4.090 ;
        RECT  4.830 0.975 6.80 1.205 ;
    END
END NA4I2X4

MACRO NA4I2X2
    CLASS CORE ;
    FOREIGN NA4I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.935 4.935 3.240 ;
        END
    END BN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.395 ;
        RECT  3.870 3.160 4.210 4.080 ;
        RECT  3.890 1.640 4.285 2.020 ;
        RECT  3.540 1.640 4.285 1.870 ;
        RECT  3.540 1.110 3.880 1.870 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.055 5.725 2.630 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.240 0.520 2.850 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.835 1.620 1.175 2.395 ;
        RECT  0.745 1.620 1.175 2.025 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.685 3.795 6.030 5.280 ;
        RECT  4.630 3.740 4.975 5.280 ;
        RECT  3.145 3.730 3.500 5.280 ;
        RECT  1.460 3.135 1.800 5.280 ;
        RECT  0.195 3.890 0.540 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.935 -0.400 6.275 0.710 ;
        RECT  4.290 -0.400 4.635 0.970 ;
        RECT  2.750 -0.400 3.090 1.330 ;
        RECT  1.270 -0.400 1.610 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.105 1.635 1.335 ;
        RECT  0.180 1.105 0.530 1.455 ;
        RECT  1.405 1.655 1.910 2.010 ;
        RECT  1.405 1.105 1.635 2.905 ;
        RECT  0.850 2.675 1.635 2.905 ;
        RECT  0.850 2.675 1.080 3.460 ;
        RECT  0.735 3.105 1.080 3.460 ;
        RECT  2.030 0.865 2.450 1.205 ;
        RECT  2.220 0.865 2.450 2.690 ;
        RECT  2.220 2.445 3.825 2.690 ;
        RECT  2.605 2.445 3.825 2.785 ;
        RECT  2.605 2.445 2.955 3.365 ;
        RECT  4.940 1.365 5.280 1.705 ;
        RECT  4.940 1.475 6.185 1.705 ;
        RECT  5.955 2.175 6.355 2.515 ;
        RECT  5.955 1.475 6.185 3.235 ;
        RECT  5.620 2.895 6.185 3.235 ;
        RECT  4.865 0.630 5.705 0.915 ;
        RECT  5.475 0.630 5.705 1.170 ;
        RECT  5.475 0.940 6.645 1.170 ;
        RECT  6.415 0.940 6.645 1.700 ;
        RECT  6.585 1.345 6.815 4.135 ;
        RECT  6.410 3.790 6.815 4.135 ;
    END
END NA4I2X2

MACRO NA4I2X1
    CLASS CORE ;
    FOREIGN NA4I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.680 0.935 2.025 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.255 1.455 2.670 ;
        END
    END D
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.930 1.920 4.295 3.240 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.885 4.975 2.655 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.772  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.125 2.930 3.700 3.160 ;
        RECT  3.470 1.640 3.700 3.160 ;
        RECT  2.875 1.640 3.700 2.020 ;
        RECT  3.125 2.930 3.465 3.800 ;
        RECT  2.875 1.530 3.215 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.055 3.800 5.400 5.280 ;
        RECT  3.885 3.900 4.230 5.280 ;
        RECT  1.595 3.900 1.935 5.280 ;
        RECT  0.275 3.700 0.615 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.165 -0.400 5.450 0.710 ;
        RECT  3.635 -0.400 3.965 0.970 ;
        RECT  1.505 -0.400 1.845 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.515 1.110 0.855 1.450 ;
        RECT  0.515 1.205 1.960 1.450 ;
        RECT  1.730 1.855 2.180 2.195 ;
        RECT  1.730 1.205 1.960 3.170 ;
        RECT  0.835 2.940 1.960 3.170 ;
        RECT  0.835 2.940 1.175 3.280 ;
        RECT  2.305 0.630 2.645 0.960 ;
        RECT  2.410 0.630 2.645 4.240 ;
        RECT  2.410 2.360 3.240 2.700 ;
        RECT  2.410 2.360 2.680 4.240 ;
        RECT  2.410 3.900 2.750 4.240 ;
        RECT  4.235 1.305 4.545 1.630 ;
        RECT  4.235 1.325 4.575 1.630 ;
        RECT  4.235 1.400 5.465 1.630 ;
        RECT  5.235 2.205 5.650 2.545 ;
        RECT  5.235 1.400 5.465 3.220 ;
        RECT  5.045 2.880 5.465 3.220 ;
        RECT  4.195 0.630 4.935 0.915 ;
        RECT  4.705 0.630 4.935 1.135 ;
        RECT  4.745 0.940 6.130 1.170 ;
        RECT  5.780 0.940 6.130 1.360 ;
        RECT  5.900 0.940 6.130 4.185 ;
        RECT  5.780 3.840 6.130 4.185 ;
    END
END NA4I2X1

MACRO NA4I2X0
    CLASS CORE ;
    FOREIGN NA4I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.690 0.520 2.300 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.599  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.655 2.020 ;
        RECT  3.110 3.630 3.505 3.960 ;
        RECT  3.275 1.330 3.505 3.960 ;
        RECT  2.815 1.330 3.505 1.670 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.415 2.670 ;
        END
    END D
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.875 2.090 4.305 2.650 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.360 4.975 3.240 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 3.440 6.120 5.280 ;
        RECT  3.740 2.880 4.080 5.280 ;
        RECT  1.580 3.530 1.920 5.280 ;
        RECT  0.180 2.875 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.100 -0.400 5.440 0.710 ;
        RECT  3.615 -0.400 3.960 0.970 ;
        RECT  2.815 -0.400 3.155 0.970 ;
        RECT  1.210 -0.400 1.550 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.520 1.460 ;
        RECT  0.180 1.225 2.015 1.460 ;
        RECT  1.645 1.225 2.015 1.565 ;
        RECT  1.645 1.225 1.875 3.165 ;
        RECT  0.880 2.935 1.875 3.165 ;
        RECT  0.880 2.935 1.110 3.760 ;
        RECT  0.880 3.420 1.220 3.760 ;
        RECT  2.015 0.630 2.475 0.970 ;
        RECT  2.245 2.360 3.045 2.700 ;
        RECT  2.245 0.630 2.475 3.870 ;
        RECT  2.245 3.530 2.735 3.870 ;
        RECT  4.175 1.370 4.525 1.670 ;
        RECT  4.175 1.385 4.555 1.670 ;
        RECT  4.175 1.400 5.435 1.670 ;
        RECT  5.205 1.760 5.645 2.100 ;
        RECT  5.205 1.400 5.435 3.870 ;
        RECT  4.770 3.530 5.435 3.870 ;
        RECT  4.190 0.630 4.870 0.915 ;
        RECT  4.640 0.630 4.870 1.170 ;
        RECT  4.640 0.940 6.045 1.170 ;
        RECT  5.690 0.940 6.045 1.455 ;
        RECT  5.715 1.240 6.105 1.470 ;
        RECT  5.875 1.240 6.105 2.980 ;
        RECT  5.665 2.640 6.105 2.980 ;
    END
END NA4I2X0

MACRO NA4I1X4
    CLASS CORE ;
    FOREIGN NA4I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.319  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.575 2.290 6.915 2.660 ;
        RECT  6.425 2.830 6.830 3.240 ;
        RECT  6.575 2.290 6.830 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.640 0.575 2.095 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.870  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.390 3.050 6.195 3.390 ;
        RECT  5.965 1.630 6.195 3.390 ;
        RECT  5.395 1.630 6.195 2.020 ;
        RECT  5.395 1.435 5.740 2.020 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.210 3.460 8.705 3.955 ;
        END
    END AN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.325 1.460 2.710 ;
        RECT  0.755 2.240 1.165 2.710 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  6.420 4.170 7.880 5.280 ;
        RECT  5.020 3.730 5.385 5.280 ;
        RECT  3.775 3.695 4.115 5.280 ;
        RECT  0.315 4.165 1.775 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.035 -0.400 8.375 0.715 ;
        RECT  6.145 -0.400 6.485 0.710 ;
        RECT  4.365 -0.400 4.705 1.180 ;
        RECT  1.375 -0.400 2.865 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.075 1.680 1.410 ;
        RECT  1.450 1.075 1.680 1.990 ;
        RECT  1.450 1.760 2.245 1.990 ;
        RECT  1.785 1.760 2.245 2.235 ;
        RECT  3.290 2.330 3.875 2.670 ;
        RECT  0.875 2.960 2.245 3.190 ;
        RECT  0.875 2.960 1.215 3.770 ;
        RECT  2.015 1.760 2.245 4.250 ;
        RECT  3.290 2.330 3.545 4.250 ;
        RECT  2.015 4.020 3.545 4.250 ;
        RECT  1.980 1.185 2.865 1.525 ;
        RECT  2.625 1.185 2.865 3.790 ;
        RECT  3.295 1.280 3.640 2.100 ;
        RECT  2.625 1.800 3.640 2.100 ;
        RECT  2.625 1.870 4.965 2.100 ;
        RECT  4.730 1.870 4.965 2.650 ;
        RECT  4.730 2.310 5.735 2.650 ;
        RECT  2.625 1.800 2.990 3.790 ;
        RECT  3.095 0.630 4.105 0.915 ;
        RECT  4.935 0.975 7.675 1.205 ;
        RECT  7.150 0.975 7.675 1.315 ;
        RECT  3.875 0.630 4.105 1.640 ;
        RECT  4.935 0.975 5.165 1.640 ;
        RECT  3.875 1.410 5.165 1.640 ;
        RECT  7.150 0.975 7.380 3.760 ;
        RECT  6.980 3.420 7.380 3.760 ;
        RECT  8.030 1.170 8.375 1.515 ;
        RECT  7.610 1.865 8.260 2.210 ;
        RECT  8.030 1.170 8.260 3.220 ;
        RECT  8.025 1.865 8.260 3.220 ;
        RECT  8.025 2.880 8.645 3.220 ;
        RECT  2.625 1.870 3.40 2.100 ;
        RECT  4.935 0.975 6.90 1.205 ;
    END
END NA4I1X4

MACRO NA4I1X2
    CLASS CORE ;
    FOREIGN NA4I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.090 1.630 1.380 2.340 ;
        RECT  0.755 1.630 1.380 2.020 ;
        END
    END D
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.345 3.475 6.815 4.010 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.240 0.685 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.163  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.955 4.865 3.250 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 1.640 4.285 3.360 ;
        RECT  3.765 3.125 4.105 4.045 ;
        RECT  3.905 1.640 4.285 2.020 ;
        RECT  3.560 1.640 4.285 1.870 ;
        RECT  3.560 1.150 3.900 1.870 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.525 3.730 5.995 5.280 ;
        RECT  3.005 4.065 3.345 5.280 ;
        RECT  0.180 3.635 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.605 -0.400 5.950 0.955 ;
        RECT  4.310 -0.400 4.660 1.035 ;
        RECT  2.790 -0.400 3.130 1.220 ;
        RECT  1.270 -0.400 1.610 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.095 1.840 1.325 ;
        RECT  0.180 1.095 0.525 1.435 ;
        RECT  1.610 1.480 2.080 1.825 ;
        RECT  1.610 1.095 1.840 3.235 ;
        RECT  0.740 2.860 1.840 3.235 ;
        RECT  2.070 0.800 2.555 1.140 ;
        RECT  2.325 0.800 2.555 2.700 ;
        RECT  2.490 2.455 3.825 2.795 ;
        RECT  2.490 2.455 2.830 3.675 ;
        RECT  4.890 0.630 5.355 0.915 ;
        RECT  5.095 0.630 5.355 1.775 ;
        RECT  5.095 1.435 5.980 1.775 ;
        RECT  5.095 0.630 5.325 3.295 ;
        RECT  5.095 2.935 5.425 3.295 ;
        RECT  6.395 0.720 6.750 1.060 ;
        RECT  6.395 0.720 6.635 2.495 ;
        RECT  5.555 2.155 6.635 2.495 ;
        RECT  6.405 0.720 6.635 3.245 ;
        RECT  6.405 2.905 6.750 3.245 ;
    END
END NA4I1X2

MACRO NA4I1X1
    CLASS CORE ;
    FOREIGN NA4I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.163  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.090 1.620 1.375 2.210 ;
        RECT  0.755 1.620 1.375 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.163  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.250 0.740 2.640 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.740 2.300 6.185 2.755 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.955 4.235 3.240 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.775  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.425 1.640 3.655 3.180 ;
        RECT  3.125 2.930 3.465 3.815 ;
        RECT  2.845 1.640 3.655 2.020 ;
        RECT  2.845 1.480 3.195 2.020 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.210 3.760 5.555 5.280 ;
        RECT  3.885 3.715 4.230 5.280 ;
        RECT  1.595 3.900 1.935 5.280 ;
        RECT  0.270 3.700 0.610 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.955 -0.400 5.300 0.970 ;
        RECT  3.600 -0.400 3.950 0.970 ;
        RECT  2.870 -0.400 3.210 0.970 ;
        RECT  1.270 -0.400 1.610 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.095 1.835 1.380 ;
        RECT  0.180 1.095 0.520 1.435 ;
        RECT  1.605 1.260 2.035 1.600 ;
        RECT  1.605 1.095 1.835 3.265 ;
        RECT  0.835 2.925 1.835 3.265 ;
        RECT  2.070 0.630 2.530 0.970 ;
        RECT  2.300 0.630 2.530 4.240 ;
        RECT  2.300 2.360 3.195 2.700 ;
        RECT  2.300 2.360 2.565 4.240 ;
        RECT  2.300 3.900 2.750 4.240 ;
        RECT  4.180 0.630 4.725 0.915 ;
        RECT  4.465 0.630 4.725 1.625 ;
        RECT  4.465 1.330 5.295 1.625 ;
        RECT  4.465 0.630 4.695 3.290 ;
        RECT  4.465 2.950 4.785 3.290 ;
        RECT  5.780 0.720 6.120 1.060 ;
        RECT  5.385 1.840 6.010 2.070 ;
        RECT  5.780 0.720 6.010 2.070 ;
        RECT  4.930 2.010 5.510 2.350 ;
        RECT  5.280 1.855 5.510 3.270 ;
        RECT  5.280 2.985 6.110 3.270 ;
    END
END NA4I1X1

MACRO NA4I1X0
    CLASS CORE ;
    FOREIGN NA4I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.690 0.515 2.300 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.589  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.635 2.000 ;
        RECT  3.275 1.640 3.605 2.020 ;
        RECT  3.275 1.330 3.505 2.770 ;
        RECT  3.110 3.530 3.450 3.870 ;
        RECT  3.250 2.635 3.480 3.815 ;
        RECT  2.815 1.330 3.505 1.670 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.415 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.830 2.125 4.235 2.650 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.570 2.275 6.175 2.590 ;
        RECT  5.595 2.170 6.175 2.590 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.085 3.420 5.425 5.280 ;
        RECT  3.710 2.880 4.050 5.280 ;
        RECT  1.580 3.530 1.920 5.280 ;
        RECT  0.180 2.875 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.345 -0.400 5.685 0.710 ;
        RECT  3.615 -0.400 3.955 0.970 ;
        RECT  2.815 -0.400 3.155 0.970 ;
        RECT  1.210 -0.400 1.550 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.520 1.460 ;
        RECT  0.180 1.225 2.015 1.460 ;
        RECT  1.730 1.150 2.015 1.490 ;
        RECT  1.645 1.225 1.875 3.165 ;
        RECT  0.880 2.935 1.875 3.165 ;
        RECT  0.880 2.935 1.110 3.760 ;
        RECT  0.880 3.420 1.220 3.760 ;
        RECT  2.015 0.630 2.475 0.920 ;
        RECT  2.245 2.175 3.045 2.515 ;
        RECT  2.245 0.630 2.475 3.870 ;
        RECT  2.245 3.530 2.735 3.870 ;
        RECT  4.185 0.630 4.525 1.500 ;
        RECT  4.465 1.265 4.945 1.575 ;
        RECT  4.465 1.265 4.930 1.605 ;
        RECT  4.465 1.265 4.695 3.760 ;
        RECT  4.385 3.420 4.725 3.760 ;
        RECT  5.145 1.690 5.685 1.920 ;
        RECT  5.345 1.170 5.685 1.920 ;
        RECT  4.925 1.840 5.365 2.170 ;
        RECT  4.925 1.840 5.210 2.210 ;
        RECT  4.925 1.840 5.155 3.110 ;
        RECT  5.710 2.820 6.050 3.110 ;
        RECT  4.925 2.825 6.050 3.110 ;
    END
END NA4I1X0

MACRO NA3X4
    CLASS CORE ;
    FOREIGN NA3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.030 0.760 2.370 ;
        RECT  0.125 1.640 0.505 2.370 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.570 2.180 7.910 2.520 ;
        RECT  7.570 0.630 7.805 2.520 ;
        RECT  5.750 0.630 7.805 0.860 ;
        RECT  3.255 2.550 6.090 2.780 ;
        RECT  5.750 0.630 6.090 2.780 ;
        RECT  3.255 0.630 3.590 2.780 ;
        RECT  1.535 0.630 3.590 0.860 ;
        RECT  1.385 1.640 1.770 2.520 ;
        RECT  1.535 0.630 1.770 2.520 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.326  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.100 2.960 8.440 3.880 ;
        RECT  0.900 3.010 8.440 3.240 ;
        RECT  6.660 2.960 8.440 3.240 ;
        RECT  6.935 1.090 7.165 3.240 ;
        RECT  6.660 2.960 7.000 3.880 ;
        RECT  6.660 1.090 7.165 1.430 ;
        RECT  5.165 3.010 5.560 3.880 ;
        RECT  3.780 3.010 4.120 3.880 ;
        RECT  2.340 2.960 2.680 3.880 ;
        RECT  2.175 1.090 2.680 1.410 ;
        RECT  2.175 1.090 2.405 3.240 ;
        RECT  0.900 2.960 2.680 3.240 ;
        RECT  0.900 2.960 1.240 3.880 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 1.640 3.025 2.675 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.820 2.960 9.160 5.280 ;
        RECT  7.380 3.470 7.720 5.280 ;
        RECT  5.940 3.470 6.280 5.280 ;
        RECT  4.500 3.470 4.840 5.280 ;
        RECT  3.060 3.470 3.400 5.280 ;
        RECT  1.620 3.470 1.960 5.280 ;
        RECT  0.180 2.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.280 -0.400 8.620 1.570 ;
        RECT  5.035 -0.400 5.420 1.875 ;
        RECT  3.955 -0.400 4.295 1.870 ;
        RECT  0.725 -0.400 1.060 1.570 ;
        RECT  0.720 -0.400 1.060 1.040 ;
        END
    END gnd!
END NA3X4

MACRO NA3X2
    CLASS CORE ;
    FOREIGN NA3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.030 0.760 2.370 ;
        RECT  0.125 1.640 0.505 2.370 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.133  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.780 2.745 4.285 3.620 ;
        RECT  0.900 2.750 4.285 2.980 ;
        RECT  2.340 2.745 2.680 3.620 ;
        RECT  2.175 1.090 2.680 1.410 ;
        RECT  2.175 1.090 2.405 2.980 ;
        RECT  0.900 2.745 1.240 3.620 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 1.640 3.025 2.315 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 0.630 3.590 2.520 ;
        RECT  1.535 0.630 3.590 0.860 ;
        RECT  1.385 1.640 1.770 2.520 ;
        RECT  1.535 0.630 1.770 2.520 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.515 2.700 4.840 5.280 ;
        RECT  3.060 3.210 3.400 5.280 ;
        RECT  1.620 3.210 1.960 5.280 ;
        RECT  0.180 2.700 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.920 -0.400 4.260 1.570 ;
        RECT  0.725 -0.400 1.060 1.570 ;
        RECT  0.720 -0.400 1.060 1.040 ;
        END
    END gnd!
END NA3X2

MACRO NA3X1
    CLASS CORE ;
    FOREIGN NA3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.575  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 3.930 2.340 4.250 ;
        RECT  2.000 2.950 2.230 4.250 ;
        RECT  1.505 1.030 2.180 1.520 ;
        RECT  1.840 0.710 2.180 1.520 ;
        RECT  0.740 2.950 2.230 3.180 ;
        RECT  1.505 1.030 1.735 3.180 ;
        RECT  1.385 1.030 2.180 1.410 ;
        RECT  0.740 2.950 1.080 3.760 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.965 1.955 2.395 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.225 1.275 2.720 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.346  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.340 0.525 2.680 ;
        RECT  0.125 2.340 0.505 3.340 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.175 4.170 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.180 -0.400 0.520 1.520 ;
        END
    END gnd!
END NA3X1

MACRO NA3X0
    CLASS CORE ;
    FOREIGN NA3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.965 1.980 2.395 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.102  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 3.810 2.340 4.150 ;
        RECT  2.000 3.160 2.230 4.150 ;
        RECT  1.505 1.170 2.180 1.510 ;
        RECT  0.735 3.160 2.230 3.390 ;
        RECT  1.385 1.030 1.765 1.410 ;
        RECT  1.505 1.030 1.735 3.390 ;
        RECT  0.735 3.160 1.040 3.500 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.225 1.245 2.725 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.640 0.525 2.980 ;
        RECT  0.125 2.640 0.505 3.340 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.455 4.170 1.640 5.280 ;
        RECT  1.300 3.810 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.180 -0.400 0.520 1.510 ;
        END
    END gnd!
END NA3X0

MACRO NA3I2X4
    CLASS CORE ;
    FOREIGN NA3I2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.590  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.995 1.135 2.640 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.452  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.875 2.010 3.200 2.345 ;
        RECT  1.875 1.665 2.365 2.345 ;
        RECT  1.875 1.640 2.345 2.345 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.590  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.935 1.995 9.500 2.640 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.135  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.395 2.920 8.075 3.260 ;
        RECT  7.725 1.510 8.065 1.850 ;
        RECT  6.215 1.510 8.065 1.770 ;
        RECT  6.395 2.860 7.465 3.260 ;
        RECT  6.395 2.860 6.735 4.140 ;
        RECT  6.215 1.385 6.720 1.770 ;
        RECT  6.215 1.385 6.450 3.095 ;
        RECT  4.960 2.865 7.465 3.095 ;
        RECT  4.955 2.910 5.295 3.250 ;
        RECT  3.885 2.930 5.295 3.160 ;
        RECT  2.075 3.035 4.040 3.265 ;
        RECT  3.820 2.980 8.075 3.095 ;
        RECT  3.515 3.035 3.855 3.365 ;
        RECT  2.075 3.035 3.855 3.320 ;
        RECT  2.075 3.035 2.415 3.385 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.435 4.160 9.900 5.280 ;
        RECT  7.115 3.650 7.455 5.280 ;
        RECT  5.675 3.325 6.015 5.280 ;
        RECT  4.235 3.620 4.575 5.280 ;
        RECT  2.795 3.585 3.135 5.280 ;
        RECT  0.180 4.160 1.655 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.435 -0.400 9.890 0.710 ;
        RECT  2.895 -0.400 3.185 1.040 ;
        RECT  2.865 -0.400 3.185 1.010 ;
        RECT  0.195 -0.400 1.700 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.560 0.630 5.270 0.860 ;
        RECT  2.115 0.830 2.475 1.410 ;
        RECT  4.930 0.630 5.270 1.200 ;
        RECT  2.115 1.220 2.745 1.410 ;
        RECT  2.115 1.180 2.710 1.410 ;
        RECT  2.530 1.270 3.900 1.500 ;
        RECT  3.560 0.630 3.900 1.670 ;
        RECT  0.795 1.220 1.135 1.575 ;
        RECT  0.795 1.335 1.605 1.575 ;
        RECT  1.365 1.335 1.605 2.805 ;
        RECT  3.435 2.290 5.510 2.630 ;
        RECT  1.365 2.575 3.665 2.805 ;
        RECT  1.365 1.335 1.595 3.100 ;
        RECT  0.745 2.870 1.595 3.100 ;
        RECT  0.745 2.870 1.085 3.760 ;
        RECT  5.650 0.635 7.440 0.900 ;
        RECT  5.650 0.635 5.990 1.045 ;
        RECT  7.100 0.635 7.440 1.240 ;
        RECT  4.270 1.455 5.985 1.795 ;
        RECT  5.650 0.635 5.985 1.880 ;
        RECT  8.995 1.220 9.335 1.575 ;
        RECT  8.465 1.335 9.335 1.575 ;
        RECT  8.465 1.335 8.705 2.455 ;
        RECT  6.680 2.115 8.705 2.455 ;
        RECT  8.475 1.335 8.705 3.100 ;
        RECT  8.475 2.870 9.335 3.100 ;
        RECT  8.995 2.870 9.335 3.760 ;
        RECT  3.435 2.290 4.50 2.630 ;
        RECT  1.365 2.575 2.60 2.805 ;
        RECT  6.680 2.115 7.80 2.455 ;
    END
END NA3I2X4

MACRO NA3I2X2
    CLASS CORE ;
    FOREIGN NA3I2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.300  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.420 0.520 2.045 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.704  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.675 1.740 5.015 2.190 ;
        RECT  4.100 1.740 5.015 1.970 ;
        RECT  4.100 0.630 4.330 1.970 ;
        RECT  2.160 0.630 4.330 0.860 ;
        RECT  1.400 1.805 2.395 2.035 ;
        RECT  2.160 0.630 2.395 2.035 ;
        RECT  2.015 1.640 2.395 2.035 ;
        RECT  1.400 1.805 1.745 2.125 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.141  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.440 2.880 4.780 3.740 ;
        RECT  2.980 2.880 4.780 3.115 ;
        RECT  1.540 2.815 3.665 3.055 ;
        RECT  3.435 1.630 3.665 3.115 ;
        RECT  3.265 1.090 3.495 2.020 ;
        RECT  2.980 2.815 3.320 3.740 ;
        RECT  2.975 1.090 3.495 1.400 ;
        RECT  1.540 2.815 1.880 3.740 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.720 1.635 6.175 2.170 ;
        END
    END BN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.200 4.135 5.540 5.280 ;
        RECT  3.720 3.345 4.060 5.280 ;
        RECT  2.260 3.285 2.615 5.280 ;
        RECT  0.780 4.140 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.560 -0.400 4.900 1.510 ;
        RECT  1.400 -0.400 1.745 1.565 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.640 0.805 0.980 1.150 ;
        RECT  0.750 0.805 0.980 2.585 ;
        RECT  2.855 2.250 3.205 2.585 ;
        RECT  0.220 2.355 3.205 2.585 ;
        RECT  0.220 2.355 0.580 3.740 ;
        RECT  5.245 0.830 5.795 1.170 ;
        RECT  3.955 2.200 4.295 2.650 ;
        RECT  3.955 2.420 5.475 2.650 ;
        RECT  5.245 0.830 5.475 3.050 ;
        RECT  5.245 2.820 6.105 3.050 ;
        RECT  5.760 2.820 6.105 3.735 ;
        RECT  0.220 2.355 2.50 2.585 ;
    END
END NA3I2X2

MACRO NA3I2X1
    CLASS CORE ;
    FOREIGN NA3I2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.600 2.855 3.185 3.270 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.225 1.565 3.700 2.070 ;
        RECT  3.225 1.545 3.670 2.070 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.955 0.455 3.240 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.294  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.685 2.855 2.370 3.240 ;
        RECT  0.685 1.360 2.115 1.675 ;
        RECT  0.685 1.360 1.135 2.035 ;
        RECT  0.685 1.360 0.915 3.240 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.330 4.075 3.675 5.280 ;
        RECT  0.185 4.170 1.590 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.215 -0.400 3.560 0.720 ;
        RECT  0.185 -0.400 0.535 1.170 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.420 0.720 2.760 2.165 ;
        RECT  1.790 1.905 2.760 2.165 ;
        RECT  2.560 3.545 2.910 4.230 ;
        RECT  1.820 3.890 2.910 4.230 ;
        RECT  3.900 1.120 4.230 1.450 ;
        RECT  1.145 2.270 1.430 2.625 ;
        RECT  1.145 2.395 4.230 2.625 ;
        RECT  3.945 1.120 4.230 3.655 ;
        RECT  3.890 2.395 4.230 3.655 ;
        RECT  1.145 2.395 3.70 2.625 ;
    END
END NA3I2X1

MACRO NA3I2X0
    CLASS CORE ;
    FOREIGN NA3I2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.250 3.065 2.640 ;
        RECT  2.685 1.840 3.065 2.640 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.035  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.690 3.435 2.395 3.910 ;
        RECT  1.355 1.170 1.980 1.460 ;
        RECT  1.690 3.130 1.920 3.910 ;
        RECT  1.345 3.130 1.920 3.360 ;
        RECT  1.345 2.820 1.585 3.360 ;
        RECT  1.355 1.170 1.585 3.360 ;
        RECT  0.455 2.820 1.585 3.050 ;
        RECT  0.455 2.820 0.795 3.160 ;
        END
    END Q
    PIN BN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.355 1.690 3.695 2.030 ;
        RECT  3.275 3.440 3.655 3.910 ;
        RECT  3.275 2.945 3.525 3.910 ;
        RECT  3.295 1.800 3.525 3.910 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.600 2.345 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.585 -0.400 3.925 0.710 ;
        RECT  0.190 -0.400 0.530 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.205 4.140 3.545 5.280 ;
        RECT  0.365 3.830 1.460 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.210 1.170 2.680 1.510 ;
        RECT  2.210 1.170 2.440 1.920 ;
        RECT  1.815 1.690 2.440 1.920 ;
        RECT  1.815 1.690 2.100 2.900 ;
        RECT  1.815 2.670 2.380 2.900 ;
        RECT  2.150 2.870 2.745 3.155 ;
        RECT  0.840 0.630 3.270 0.860 ;
        RECT  3.040 0.630 3.270 1.170 ;
        RECT  3.040 0.940 4.230 1.170 ;
        RECT  3.890 0.940 4.230 1.510 ;
        RECT  0.840 0.630 1.125 2.400 ;
        RECT  3.805 2.640 4.230 2.925 ;
        RECT  3.945 0.940 4.230 2.950 ;
        RECT  3.830 2.640 4.230 2.950 ;
        RECT  0.840 0.630 2.70 0.860 ;
    END
END NA3I2X0

MACRO NA3I1X4
    CLASS CORE ;
    FOREIGN NA3I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.380  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.875 2.010 3.295 2.345 ;
        RECT  1.875 1.640 2.395 2.345 ;
        END
    END C
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.590  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.995 1.135 2.640 ;
        END
    END AN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.242  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.765 0.700 8.010 3.330 ;
        RECT  7.040 2.860 8.010 3.330 ;
        RECT  6.330 1.360 8.010 1.700 ;
        RECT  7.670 0.700 8.010 1.700 ;
        RECT  4.955 3.100 8.010 3.330 ;
        RECT  6.300 3.100 6.640 3.445 ;
        RECT  2.075 3.330 5.295 3.560 ;
        RECT  3.515 3.330 3.855 4.180 ;
        RECT  2.075 3.035 2.420 3.560 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.380  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.120 5.440 2.410 ;
        RECT  3.895 2.120 4.340 2.450 ;
        RECT  3.895 2.120 4.245 2.590 ;
        RECT  3.895 2.120 4.240 2.640 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.020 3.650 7.360 5.280 ;
        RECT  5.580 3.765 5.920 5.280 ;
        RECT  4.235 3.790 4.575 5.280 ;
        RECT  2.795 3.820 3.135 5.280 ;
        RECT  0.180 4.160 1.655 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  2.840 -0.400 3.145 0.980 ;
        RECT  2.805 -0.400 3.145 0.965 ;
        RECT  0.195 -0.400 1.665 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.525 0.730 5.220 1.100 ;
        RECT  2.080 0.825 2.440 1.410 ;
        RECT  2.080 1.180 2.715 1.410 ;
        RECT  2.530 1.210 3.865 1.440 ;
        RECT  3.525 0.730 3.865 1.650 ;
        RECT  5.600 0.770 7.290 1.110 ;
        RECT  5.600 0.770 5.940 1.695 ;
        RECT  4.235 1.355 5.940 1.695 ;
        RECT  0.760 1.220 1.605 1.575 ;
        RECT  6.090 2.200 7.500 2.545 ;
        RECT  1.365 1.220 1.605 2.805 ;
        RECT  1.365 2.575 3.665 2.805 ;
        RECT  3.435 2.575 3.665 3.100 ;
        RECT  4.470 2.640 6.325 2.870 ;
        RECT  6.090 2.200 6.325 2.870 ;
        RECT  1.365 1.220 1.595 3.100 ;
        RECT  0.745 2.870 1.595 3.100 ;
        RECT  3.435 2.870 4.700 3.100 ;
        RECT  0.745 2.870 1.085 3.760 ;
        RECT  1.365 2.575 2.30 2.805 ;
    END
END NA3I1X4

MACRO NA3I1X2
    CLASS CORE ;
    FOREIGN NA3I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.300  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.420 0.520 2.045 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.704  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.655 1.740 4.995 2.090 ;
        RECT  4.100 1.740 4.995 1.970 ;
        RECT  4.100 0.630 4.330 1.970 ;
        RECT  2.160 0.630 4.330 0.860 ;
        RECT  1.400 1.805 2.395 2.035 ;
        RECT  2.160 0.630 2.395 2.035 ;
        RECT  2.015 1.640 2.395 2.035 ;
        RECT  1.400 1.805 1.745 2.125 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.141  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.420 2.880 4.760 3.740 ;
        RECT  2.980 2.880 4.760 3.110 ;
        RECT  1.540 2.815 3.665 3.055 ;
        RECT  3.435 1.630 3.665 3.110 ;
        RECT  3.265 1.090 3.495 2.020 ;
        RECT  2.980 2.815 3.320 3.740 ;
        RECT  2.975 1.090 3.495 1.400 ;
        RECT  1.540 2.815 1.880 3.740 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.704  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.200 4.445 2.650 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.140 2.815 5.480 5.280 ;
        RECT  3.700 3.345 4.040 5.280 ;
        RECT  2.260 3.285 2.615 5.280 ;
        RECT  0.780 4.140 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.560 -0.400 4.900 1.510 ;
        RECT  1.400 -0.400 1.745 1.565 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.640 0.805 0.980 1.150 ;
        RECT  0.750 0.805 0.980 2.585 ;
        RECT  2.855 2.250 3.205 2.585 ;
        RECT  0.220 2.355 3.205 2.585 ;
        RECT  0.220 2.355 0.580 3.740 ;
        RECT  0.220 2.355 2.20 2.585 ;
    END
END NA3I1X2

MACRO NA3I1X1
    CLASS CORE ;
    FOREIGN NA3I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.980 1.635 3.655 2.070 ;
        END
    END AN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.352  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.605 0.455 2.325 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.352  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.145 2.180 1.765 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.481  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.685 1.380 2.140 1.720 ;
        RECT  1.795 0.700 2.140 1.720 ;
        RECT  1.685 2.860 2.040 3.740 ;
        RECT  0.180 2.860 2.040 3.240 ;
        RECT  0.180 2.810 0.915 3.240 ;
        RECT  0.685 1.380 0.915 3.240 ;
        RECT  0.180 2.810 0.520 3.740 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.460 2.815 2.800 5.280 ;
        RECT  0.940 3.470 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.190 -0.400 3.535 0.820 ;
        RECT  0.180 -0.400 0.520 1.185 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.500 1.110 2.840 1.450 ;
        RECT  2.500 1.110 2.750 2.530 ;
        RECT  2.180 2.190 2.750 2.530 ;
        RECT  2.180 2.300 3.565 2.530 ;
        RECT  3.220 2.300 3.565 3.180 ;
    END
END NA3I1X1

MACRO NA3I1X0
    CLASS CORE ;
    FOREIGN NA3I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.615 0.455 2.315 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.145 2.180 1.765 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.108  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.685 1.105 1.940 1.445 ;
        RECT  0.180 3.490 1.840 3.855 ;
        RECT  0.685 3.470 1.840 3.855 ;
        RECT  0.685 1.105 0.915 3.855 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.575 2.655 ;
        RECT  2.290 1.885 2.575 2.655 ;
        END
    END AN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.170 2.985 2.510 3.325 ;
        RECT  2.170 2.985 2.400 5.280 ;
        RECT  0.830 4.170 1.170 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 0.710 ;
        RECT  0.180 -0.400 0.535 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.375 0.630 2.400 0.875 ;
        RECT  2.170 0.630 2.400 1.170 ;
        RECT  2.170 0.940 3.035 1.170 ;
        RECT  2.630 0.940 3.035 1.510 ;
        RECT  2.805 0.940 3.035 4.170 ;
        RECT  2.630 3.830 3.035 4.170 ;
    END
END NA3I1X0

MACRO NA2X4
    CLASS CORE ;
    FOREIGN NA2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.024  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.060 1.950 5.400 3.580 ;
        RECT  0.740 1.950 5.400 2.235 ;
        RECT  3.910 1.240 4.250 2.235 ;
        RECT  3.610 1.950 3.970 3.580 ;
        RECT  2.180 1.950 2.520 3.580 ;
        RECT  1.385 1.240 1.950 2.235 ;
        RECT  0.740 1.950 1.080 3.580 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.900 0.510 2.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.785 1.640 6.175 2.410 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.770 2.640 6.120 5.280 ;
        RECT  4.325 2.660 4.695 5.280 ;
        RECT  2.900 2.660 3.240 5.280 ;
        RECT  1.460 2.660 1.800 5.280 ;
        RECT  0.180 3.980 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.100 -0.400 5.440 1.720 ;
        RECT  2.760 -0.400 3.100 1.580 ;
        RECT  0.420 -0.400 0.760 1.670 ;
        END
    END gnd!
END NA2X4

MACRO NA2X2
    CLASS CORE ;
    FOREIGN NA2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.705 2.860 3.935 ;
        RECT  2.630 2.260 2.860 3.935 ;
        RECT  2.290 2.260 2.860 2.600 ;
        RECT  0.115 1.630 0.560 2.030 ;
        RECT  0.115 1.630 0.345 3.935 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.175 1.305 2.695 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.512  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 3.135 2.400 3.475 ;
        RECT  1.535 1.030 1.765 3.475 ;
        RECT  1.330 1.030 1.765 1.510 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.180 4.170 2.960 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.560 -0.400 2.900 1.510 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
END NA2X2

MACRO NA2X1
    CLASS CORE ;
    FOREIGN NA2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.630 0.545 2.015 ;
        RECT  0.115 1.630 0.525 2.215 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.110 1.305 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.924  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.780 2.860 1.765 3.200 ;
        RECT  1.535 1.030 1.765 3.200 ;
        RECT  1.330 1.030 1.765 1.510 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  0.180 4.170 1.710 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
END NA2X1

MACRO NA2X0
    CLASS CORE ;
    FOREIGN NA2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.565 0.525 3.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.220 1.225 2.740 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.518  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.330 1.030 1.765 1.410 ;
        RECT  0.780 3.090 1.685 3.430 ;
        RECT  1.455 1.030 1.685 3.430 ;
        RECT  1.330 1.030 1.685 1.510 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  1.370 3.890 1.710 5.280 ;
        RECT  0.180 3.835 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  0.180 -0.400 0.520 0.930 ;
        END
    END gnd!
END NA2X0

MACRO NA2I1X4
    CLASS CORE ;
    FOREIGN NA2I1X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.590  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.995 1.135 2.640 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.296  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.845 3.375 2.170 ;
        RECT  1.995 1.655 2.380 2.170 ;
        RECT  1.995 1.640 2.345 2.170 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.258  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.600 1.710 6.120 1.940 ;
        RECT  5.780 0.700 6.120 1.940 ;
        RECT  4.955 2.640 5.295 3.910 ;
        RECT  5.040 1.710 5.295 3.910 ;
        RECT  2.075 2.860 5.295 3.095 ;
        RECT  4.600 1.090 4.830 1.940 ;
        RECT  4.330 1.090 4.830 1.430 ;
        RECT  3.515 2.860 3.855 3.910 ;
        RECT  3.270 2.860 3.855 3.245 ;
        RECT  2.075 2.860 3.855 3.145 ;
        RECT  2.075 2.860 2.415 3.910 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.675 2.640 6.015 5.280 ;
        RECT  4.235 3.325 4.575 5.280 ;
        RECT  2.795 3.480 3.135 5.280 ;
        RECT  0.180 3.960 1.655 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  2.955 -0.400 3.245 1.040 ;
        RECT  2.925 -0.400 3.245 1.010 ;
        RECT  0.255 -0.400 1.755 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.855 1.220 1.195 1.575 ;
        RECT  0.855 1.335 1.605 1.575 ;
        RECT  1.365 1.335 1.605 2.630 ;
        RECT  3.995 2.170 4.805 2.460 ;
        RECT  3.995 2.120 4.335 2.630 ;
        RECT  1.365 2.400 4.335 2.630 ;
        RECT  1.365 1.335 1.595 3.210 ;
        RECT  0.745 2.980 1.595 3.210 ;
        RECT  0.745 2.980 1.085 3.330 ;
        RECT  3.620 0.630 5.400 0.860 ;
        RECT  2.175 1.070 2.535 1.410 ;
        RECT  2.175 1.220 2.805 1.410 ;
        RECT  2.175 1.180 2.770 1.410 ;
        RECT  5.060 0.630 5.400 1.480 ;
        RECT  2.575 1.300 3.960 1.530 ;
        RECT  3.620 0.630 3.960 1.670 ;
        RECT  1.365 2.400 3.60 2.630 ;
    END
END NA2I1X4

MACRO NA2I1X2
    CLASS CORE ;
    FOREIGN NA2I1X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.293  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.870 0.505 2.605 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.025 1.565 3.365 2.020 ;
        RECT  2.795 0.630 3.025 1.805 ;
        RECT  1.615 0.630 3.025 0.860 ;
        RECT  1.205 1.635 1.850 2.020 ;
        RECT  1.615 0.630 1.850 2.020 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.640  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.700 2.790 3.040 3.700 ;
        RECT  1.340 2.965 3.040 3.250 ;
        RECT  2.375 2.790 3.040 3.250 ;
        RECT  2.375 1.970 2.605 3.250 ;
        RECT  2.335 1.090 2.565 2.105 ;
        RECT  2.105 1.090 2.565 1.430 ;
        RECT  1.340 2.965 1.680 4.250 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.140 4.105 3.600 5.280 ;
        RECT  0.770 3.295 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.260 -0.400 3.600 1.180 ;
        RECT  0.940 -0.400 1.280 1.170 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.020 0.520 1.640 ;
        RECT  0.180 1.400 0.975 1.640 ;
        RECT  0.735 1.400 0.975 2.590 ;
        RECT  0.735 2.250 2.145 2.590 ;
        RECT  0.735 1.400 0.965 3.065 ;
        RECT  0.180 2.835 0.965 3.065 ;
        RECT  0.180 2.835 0.520 4.250 ;
    END
END NA2I1X2

MACRO NA2I1X1
    CLASS CORE ;
    FOREIGN NA2I1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.870 0.505 2.630 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.215 1.635 1.850 2.020 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.954  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.460 0.990 3.025 1.410 ;
        RECT  1.715 2.825 2.760 3.110 ;
        RECT  2.460 0.990 2.760 3.110 ;
        RECT  2.165 0.990 3.025 1.330 ;
        RECT  1.715 2.825 2.055 3.855 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.490 3.340 2.830 5.280 ;
        RECT  0.940 3.320 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  0.980 -0.400 1.320 1.170 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.940 0.520 1.640 ;
        RECT  0.180 1.400 0.975 1.640 ;
        RECT  0.735 1.400 0.975 2.590 ;
        RECT  0.735 2.250 2.230 2.590 ;
        RECT  0.735 1.400 0.965 3.090 ;
        RECT  0.180 2.860 0.965 3.090 ;
        RECT  0.180 2.860 0.520 3.300 ;
    END
END NA2I1X1

MACRO NA2I1X0
    CLASS CORE ;
    FOREIGN NA2I1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.803  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.590 3.160 2.395 3.445 ;
        RECT  2.165 1.030 2.395 3.445 ;
        RECT  2.000 1.030 2.395 1.520 ;
        END
    END Q
    PIN AN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.160 0.570 2.645 ;
        RECT  0.125 2.115 0.505 2.645 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.805 1.640 1.215 2.220 ;
        RECT  0.755 1.640 1.215 2.020 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  1.710 3.940 2.050 5.280 ;
        RECT  0.890 3.570 1.230 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.890 -0.400 1.230 0.790 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.260 ;
        RECT  0.180 1.020 1.685 1.260 ;
        RECT  1.445 1.020 1.685 2.930 ;
        RECT  1.445 2.330 1.935 2.930 ;
        RECT  0.795 2.700 1.935 2.930 ;
        RECT  0.795 2.700 1.025 3.290 ;
        RECT  0.180 3.060 1.025 3.290 ;
        RECT  0.180 3.060 0.520 3.840 ;
    END
END NA2I1X0

MACRO MU4X4
    CLASS CORE ;
    FOREIGN MU4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.835 2.025 4.290 2.630 ;
        END
    END IN0
    PIN S1
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.196  LAYER MET1  ;
        ANTENNAGATEAREA 1.962  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.115 3.470 20.035 4.050 ;
        RECT  19.115 2.450 19.345 4.050 ;
        RECT  17.390 2.450 19.345 2.680 ;
        RECT  17.390 2.340 17.675 2.680 ;
        RECT  8.855 2.580 9.195 2.920 ;
        RECT  6.940 2.580 9.195 2.810 ;
        RECT  6.940 2.580 7.280 2.920 ;
        END
    END S1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.605 1.145 18.945 1.670 ;
        RECT  15.455 1.145 18.945 1.375 ;
        RECT  16.600 3.370 17.695 3.600 ;
        RECT  8.495 3.305 16.765 3.425 ;
        RECT  11.875 3.370 17.695 3.535 ;
        RECT  15.455 1.035 16.015 1.375 ;
        RECT  13.960 1.515 15.685 1.745 ;
        RECT  15.455 1.035 15.685 1.745 ;
        RECT  12.925 2.385 14.190 2.615 ;
        RECT  13.960 0.850 14.190 2.615 ;
        RECT  13.205 0.850 14.190 1.190 ;
        RECT  12.925 1.880 13.155 2.615 ;
        RECT  10.965 1.880 13.155 2.110 ;
        RECT  11.875 3.195 12.215 3.790 ;
        RECT  11.985 1.880 12.215 3.790 ;
        RECT  11.900 2.860 12.215 3.790 ;
        RECT  8.495 3.195 12.215 3.425 ;
        RECT  10.965 1.345 11.195 2.110 ;
        RECT  9.910 1.345 11.195 1.575 ;
        RECT  10.430 1.090 10.770 1.575 ;
        RECT  10.205 2.860 10.585 3.425 ;
        RECT  7.830 1.660 10.140 1.890 ;
        RECT  9.910 1.345 10.140 1.890 ;
        RECT  8.495 3.195 9.555 3.535 ;
        RECT  7.830 1.150 8.060 1.890 ;
        RECT  7.360 1.150 8.060 1.490 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.206  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.245 0.705 2.625 ;
        END
    END S0
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.090 1.640 1.385 2.140 ;
        RECT  0.755 1.640 1.385 2.020 ;
        END
    END IN2
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.195 1.640 3.610 1.975 ;
        RECT  3.195 1.640 3.605 2.215 ;
        END
    END IN3
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.605 1.555 6.175 2.020 ;
        END
    END IN1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  19.335 -0.400 19.675 0.710 ;
        RECT  16.865 -0.400 17.755 0.915 ;
        RECT  14.525 -0.400 14.865 1.285 ;
        RECT  11.885 -0.400 12.185 1.190 ;
        RECT  8.880 -0.400 9.220 0.970 ;
        RECT  5.860 -0.400 6.200 0.655 ;
        RECT  3.475 -0.400 3.825 0.950 ;
        RECT  0.920 -0.400 1.260 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  18.545 2.910 18.885 5.280 ;
        RECT  15.765 4.225 16.105 5.280 ;
        RECT  13.340 4.225 13.680 5.280 ;
        RECT  10.520 4.225 10.860 5.280 ;
        RECT  7.400 3.610 7.685 5.280 ;
        RECT  5.770 4.130 6.110 5.280 ;
        RECT  3.225 3.360 3.565 5.280 ;
        RECT  0.900 3.315 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.700 0.520 1.620 ;
        RECT  0.180 1.180 1.845 1.410 ;
        RECT  0.180 1.180 0.525 1.620 ;
        RECT  1.615 1.870 2.505 2.210 ;
        RECT  0.180 2.855 1.845 3.085 ;
        RECT  4.575 1.940 4.915 3.130 ;
        RECT  2.755 2.900 4.915 3.130 ;
        RECT  1.615 1.180 1.845 4.085 ;
        RECT  2.755 2.900 2.985 4.085 ;
        RECT  1.615 3.855 2.985 4.085 ;
        RECT  0.180 2.855 0.520 4.180 ;
        RECT  6.660 1.345 7.000 2.350 ;
        RECT  7.260 1.825 7.600 2.350 ;
        RECT  6.475 2.120 10.710 2.350 ;
        RECT  10.370 1.805 10.710 2.350 ;
        RECT  10.480 2.340 11.755 2.570 ;
        RECT  11.470 2.340 11.755 2.680 ;
        RECT  6.475 2.120 6.710 3.440 ;
        RECT  4.085 0.630 5.530 0.860 ;
        RECT  9.450 0.630 11.655 0.860 ;
        RECT  5.300 0.630 5.530 1.115 ;
        RECT  6.790 0.690 8.565 0.920 ;
        RECT  5.300 0.885 7.020 1.115 ;
        RECT  2.120 0.980 2.465 1.415 ;
        RECT  8.310 0.690 8.565 1.430 ;
        RECT  4.085 0.630 4.315 1.410 ;
        RECT  2.120 1.180 4.315 1.410 ;
        RECT  2.120 1.180 2.965 1.415 ;
        RECT  11.425 0.630 11.655 1.650 ;
        RECT  9.450 0.630 9.680 1.430 ;
        RECT  8.310 1.200 9.680 1.430 ;
        RECT  11.425 1.420 13.725 1.650 ;
        RECT  13.385 1.420 13.725 2.155 ;
        RECT  2.735 1.180 2.965 2.670 ;
        RECT  2.075 2.440 2.965 2.670 ;
        RECT  2.075 2.440 2.415 3.625 ;
        RECT  4.670 1.090 5.060 1.575 ;
        RECT  4.670 1.345 5.375 1.575 ;
        RECT  16.605 2.065 17.160 2.350 ;
        RECT  16.930 2.065 17.160 3.140 ;
        RECT  16.930 2.910 18.155 3.140 ;
        RECT  6.940 3.150 8.180 3.380 ;
        RECT  5.145 1.345 5.375 3.900 ;
        RECT  4.580 3.360 5.375 3.900 ;
        RECT  5.920 2.340 6.245 3.900 ;
        RECT  7.950 3.150 8.180 3.995 ;
        RECT  6.940 3.150 7.170 3.900 ;
        RECT  4.580 3.670 7.170 3.900 ;
        RECT  7.950 3.765 11.320 3.995 ;
        RECT  12.880 3.765 16.435 3.995 ;
        RECT  11.090 3.765 11.320 4.250 ;
        RECT  17.925 2.910 18.155 4.060 ;
        RECT  16.270 3.830 18.155 4.060 ;
        RECT  4.580 3.360 4.920 4.175 ;
        RECT  12.880 3.765 13.110 4.250 ;
        RECT  11.090 4.020 13.110 4.250 ;
        RECT  15.915 1.605 18.375 1.835 ;
        RECT  18.145 1.605 18.375 2.130 ;
        RECT  18.145 1.900 19.915 2.130 ;
        RECT  19.375 1.090 19.715 2.220 ;
        RECT  18.610 1.900 19.915 2.220 ;
        RECT  15.915 1.605 16.255 2.680 ;
        RECT  14.510 2.340 16.255 2.680 ;
        RECT  12.445 2.340 12.695 3.075 ;
        RECT  14.510 2.340 14.740 3.075 ;
        RECT  12.445 2.845 14.740 3.075 ;
        RECT  19.575 1.900 19.915 3.240 ;
        RECT  2.755 2.900 3.80 3.130 ;
        RECT  6.475 2.120 9.90 2.350 ;
        RECT  9.450 0.630 10.50 0.860 ;
        RECT  2.120 1.180 3.60 1.410 ;
        RECT  11.425 1.420 12.70 1.650 ;
        RECT  4.580 3.670 6.60 3.900 ;
        RECT  7.950 3.765 10.90 3.995 ;
        RECT  12.880 3.765 15.70 3.995 ;
        RECT  11.090 4.020 12.60 4.250 ;
        RECT  15.915 1.605 17.70 1.835 ;
        RECT  12.445 2.845 13.60 3.075 ;
    END
END MU4X4

MACRO MU4X2
    CLASS CORE ;
    FOREIGN MU4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.336  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.400 3.460 9.965 3.860 ;
        RECT  9.285 1.230 9.790 1.570 ;
        RECT  9.400 3.235 9.745 4.140 ;
        RECT  7.970 2.315 9.515 2.545 ;
        RECT  9.285 1.230 9.515 2.545 ;
        RECT  6.470 3.235 9.745 3.465 ;
        RECT  7.970 1.615 8.200 2.545 ;
        RECT  7.395 1.615 8.200 1.845 ;
        RECT  6.470 1.575 7.560 1.805 ;
        RECT  7.060 3.235 7.405 3.585 ;
        RECT  6.980 1.090 7.320 1.805 ;
        RECT  6.470 1.575 6.700 3.465 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.054  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.435 1.640 11.855 2.220 ;
        END
    END S1
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.020 2.270 3.665 2.640 ;
        RECT  3.020 2.250 3.395 2.640 ;
        RECT  3.020 2.240 3.380 2.640 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.947  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.250 0.660 2.625 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.505 1.615 6.175 2.035 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.000 1.625 1.340 2.205 ;
        RECT  0.755 1.625 1.340 2.020 ;
        END
    END IN0
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.625 1.640 4.235 2.040 ;
        END
    END IN2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.685 2.935 11.070 5.280 ;
        RECT  8.255 3.695 8.595 5.280 ;
        RECT  5.730 2.910 6.085 5.280 ;
        RECT  3.320 3.330 3.660 5.280 ;
        RECT  0.935 3.315 1.275 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.640 -0.400 10.995 0.970 ;
        RECT  8.215 -0.400 8.555 0.925 ;
        RECT  5.785 -0.400 6.130 0.710 ;
        RECT  3.360 -0.400 3.710 0.950 ;
        RECT  0.940 -0.400 1.280 0.915 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.845 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  1.610 1.830 2.175 2.170 ;
        RECT  0.215 2.855 1.840 3.085 ;
        RECT  4.465 1.870 4.695 3.100 ;
        RECT  2.755 2.870 4.695 3.100 ;
        RECT  1.610 1.145 1.840 4.085 ;
        RECT  0.215 2.855 0.555 3.880 ;
        RECT  2.755 2.870 2.985 4.085 ;
        RECT  1.610 3.855 2.985 4.085 ;
        RECT  4.600 1.145 4.990 1.585 ;
        RECT  5.955 2.340 6.240 2.680 ;
        RECT  4.925 2.450 6.240 2.680 ;
        RECT  4.925 1.360 5.155 3.680 ;
        RECT  4.545 3.340 5.155 3.680 ;
        RECT  6.440 0.630 7.985 0.860 ;
        RECT  4.085 0.685 5.515 0.915 ;
        RECT  5.285 0.685 5.515 1.170 ;
        RECT  8.805 0.750 10.410 0.980 ;
        RECT  7.755 0.630 7.985 1.385 ;
        RECT  6.440 0.630 6.675 1.170 ;
        RECT  5.285 0.940 6.675 1.170 ;
        RECT  8.805 0.750 9.035 1.385 ;
        RECT  7.755 1.155 9.035 1.385 ;
        RECT  4.085 0.685 4.315 1.410 ;
        RECT  2.155 1.180 4.315 1.410 ;
        RECT  2.155 1.075 2.500 1.415 ;
        RECT  10.180 0.750 10.410 1.500 ;
        RECT  10.360 1.270 10.590 2.145 ;
        RECT  8.455 1.155 8.795 2.085 ;
        RECT  10.360 1.805 10.700 2.145 ;
        RECT  2.405 1.180 2.635 2.630 ;
        RECT  2.130 2.400 2.470 3.625 ;
        RECT  11.110 1.180 11.785 1.410 ;
        RECT  11.440 1.025 11.785 1.410 ;
        RECT  9.745 1.800 10.035 2.690 ;
        RECT  10.975 1.200 11.205 2.690 ;
        RECT  9.745 2.460 11.785 2.690 ;
        RECT  6.930 2.035 7.220 3.005 ;
        RECT  9.745 1.800 9.975 3.005 ;
        RECT  6.930 2.775 9.975 3.005 ;
        RECT  11.435 2.460 11.785 3.840 ;
        RECT  2.155 1.180 3.80 1.410 ;
        RECT  9.745 2.460 10.30 2.690 ;
        RECT  6.930 2.775 8.40 3.005 ;
    END
END MU4X2

MACRO MU4X1
    CLASS CORE ;
    FOREIGN MU4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.423  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.975 2.785 7.435 3.250 ;
        RECT  6.975 2.785 7.320 4.120 ;
        RECT  6.415 1.500 7.320 1.730 ;
        RECT  6.980 1.285 7.320 1.730 ;
        RECT  6.415 2.785 7.435 3.085 ;
        RECT  6.415 1.500 6.645 3.085 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.527  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.820 3.410 9.335 3.890 ;
        END
    END S1
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.480 2.020 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.546  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.605 0.620 2.020 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.600 1.520 6.175 2.020 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.230 1.350 2.615 ;
        RECT  1.000 2.190 1.350 2.615 ;
        END
    END IN0
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.720 1.640 4.245 2.020 ;
        RECT  3.720 1.640 4.060 2.520 ;
        END
    END IN2
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.130 -0.400 8.470 1.525 ;
        RECT  5.745 -0.400 6.090 0.710 ;
        RECT  3.410 -0.400 3.760 0.915 ;
        RECT  0.980 -0.400 1.320 0.915 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.170 2.785 8.510 5.280 ;
        RECT  5.810 2.855 6.165 5.280 ;
        RECT  3.320 3.475 3.660 5.280 ;
        RECT  0.980 3.305 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.635 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  1.610 1.930 1.955 2.270 ;
        RECT  1.610 1.145 1.840 3.250 ;
        RECT  4.465 2.095 4.695 2.990 ;
        RECT  2.795 2.760 4.695 2.990 ;
        RECT  0.185 2.845 1.840 3.075 ;
        RECT  2.795 2.760 3.025 3.250 ;
        RECT  1.610 3.020 3.025 3.250 ;
        RECT  0.185 2.845 0.545 3.515 ;
        RECT  4.690 1.110 5.030 1.810 ;
        RECT  4.925 2.280 6.185 2.625 ;
        RECT  4.925 1.585 5.155 3.505 ;
        RECT  4.520 3.220 5.155 3.505 ;
        RECT  4.085 0.630 5.515 0.860 ;
        RECT  5.285 0.630 5.515 1.170 ;
        RECT  6.440 0.825 7.845 1.055 ;
        RECT  2.185 0.980 2.550 1.375 ;
        RECT  5.285 0.940 6.675 1.170 ;
        RECT  4.085 0.630 4.315 1.375 ;
        RECT  2.185 1.145 4.315 1.375 ;
        RECT  7.615 0.825 7.845 2.095 ;
        RECT  7.615 1.810 8.265 2.095 ;
        RECT  2.185 0.980 2.415 2.790 ;
        RECT  2.170 2.450 2.510 2.790 ;
        RECT  6.875 1.960 7.160 2.555 ;
        RECT  6.875 2.325 9.270 2.555 ;
        RECT  8.930 1.285 9.270 3.075 ;
        RECT  2.185 1.145 3.60 1.375 ;
        RECT  6.875 2.325 8.70 2.555 ;
    END
END MU4X1

MACRO MU4X0
    CLASS CORE ;
    FOREIGN MU4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.830 1.640 4.285 2.530 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.480 2.060 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.405  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.605 0.670 2.020 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.450 1.640 6.175 1.995 ;
        RECT  5.450 1.640 5.735 2.105 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.240 1.380 2.580 ;
        RECT  1.000 2.165 1.380 2.580 ;
        END
    END IN0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.539  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.815 2.800 7.435 3.240 ;
        RECT  6.915 1.170 7.240 1.620 ;
        RECT  6.815 1.390 7.045 3.240 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.277  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.725 3.450 9.330 3.855 ;
        END
    END S1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.180 -0.400 8.470 1.325 ;
        RECT  5.915 -0.400 6.210 0.710 ;
        RECT  3.460 -0.400 3.820 0.915 ;
        RECT  0.980 -0.400 1.320 0.915 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.130 2.775 8.470 5.280 ;
        RECT  5.775 2.850 6.115 5.280 ;
        RECT  3.340 3.325 3.680 5.280 ;
        RECT  1.025 3.270 1.365 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.635 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  4.515 1.730 4.760 2.990 ;
        RECT  2.795 2.760 4.760 2.990 ;
        RECT  1.610 1.145 1.840 3.040 ;
        RECT  0.225 2.810 1.955 3.040 ;
        RECT  1.725 1.930 1.955 3.295 ;
        RECT  2.795 2.760 3.025 3.295 ;
        RECT  1.725 3.060 3.025 3.295 ;
        RECT  0.225 2.810 0.585 3.455 ;
        RECT  4.640 1.090 5.220 1.375 ;
        RECT  6.070 2.225 6.410 2.620 ;
        RECT  4.990 2.390 6.410 2.620 ;
        RECT  4.990 1.090 5.220 3.510 ;
        RECT  4.550 3.220 5.220 3.510 ;
        RECT  4.085 0.630 5.685 0.860 ;
        RECT  6.455 0.630 7.950 0.860 ;
        RECT  5.455 0.630 5.685 1.175 ;
        RECT  2.185 0.875 2.550 1.375 ;
        RECT  6.455 0.630 6.685 1.175 ;
        RECT  5.455 0.945 6.685 1.175 ;
        RECT  4.085 0.630 4.315 1.375 ;
        RECT  2.185 1.145 4.315 1.375 ;
        RECT  7.720 0.630 7.950 1.760 ;
        RECT  7.845 1.555 8.230 1.815 ;
        RECT  2.185 0.875 2.415 2.830 ;
        RECT  2.185 2.490 2.565 2.830 ;
        RECT  7.275 1.855 7.505 2.275 ;
        RECT  7.275 2.045 9.270 2.275 ;
        RECT  8.930 1.010 9.270 3.085 ;
        RECT  2.185 1.145 3.60 1.375 ;
    END
END MU4X0

MACRO MU4IX4
    CLASS CORE ;
    FOREIGN MU4IX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.375  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 0.700 14.365 2.025 ;
        RECT  13.970 0.700 14.310 4.130 ;
        RECT  12.650 2.640 14.310 2.870 ;
        RECT  12.650 1.180 14.365 1.520 ;
        RECT  12.650 2.640 12.990 3.755 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.435 1.640 11.880 2.185 ;
        END
    END S1
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.195 1.640 3.610 1.975 ;
        RECT  3.195 1.640 3.605 2.215 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.206  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.245 0.705 2.625 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.605 1.615 6.175 2.110 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.090 1.640 1.385 2.140 ;
        RECT  0.755 1.640 1.385 2.020 ;
        END
    END IN0
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.835 2.025 4.290 2.630 ;
        END
    END IN2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.210 4.170 13.550 5.280 ;
        RECT  12.100 4.170 12.445 5.280 ;
        RECT  10.710 3.535 11.050 5.280 ;
        RECT  8.240 3.695 8.580 5.280 ;
        RECT  5.730 2.910 6.070 5.280 ;
        RECT  3.225 3.360 3.565 5.280 ;
        RECT  0.900 3.315 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.210 -0.400 13.550 0.710 ;
        RECT  11.890 -0.400 12.230 0.710 ;
        RECT  10.610 -0.400 10.965 0.960 ;
        RECT  8.240 -0.400 8.580 0.925 ;
        RECT  5.855 -0.400 6.200 0.710 ;
        RECT  3.475 -0.400 3.825 0.950 ;
        RECT  0.920 -0.400 1.260 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.700 0.520 1.620 ;
        RECT  0.180 1.180 1.845 1.410 ;
        RECT  0.180 1.180 0.525 1.620 ;
        RECT  1.615 1.870 2.505 2.210 ;
        RECT  0.180 2.855 1.845 3.085 ;
        RECT  4.575 1.940 4.915 3.130 ;
        RECT  2.755 2.900 4.915 3.130 ;
        RECT  1.615 1.180 1.845 4.085 ;
        RECT  2.755 2.900 2.985 4.085 ;
        RECT  1.615 3.855 2.985 4.085 ;
        RECT  0.180 2.855 0.520 4.180 ;
        RECT  4.670 1.090 5.060 1.630 ;
        RECT  4.670 1.400 5.375 1.630 ;
        RECT  5.920 2.340 6.260 2.680 ;
        RECT  5.145 2.450 6.260 2.680 ;
        RECT  5.145 1.400 5.375 3.690 ;
        RECT  4.580 3.360 5.375 3.690 ;
        RECT  4.580 3.360 4.920 4.175 ;
        RECT  4.085 0.630 5.530 0.860 ;
        RECT  6.455 0.630 7.985 0.860 ;
        RECT  5.300 0.630 5.530 1.170 ;
        RECT  8.810 0.750 10.370 0.980 ;
        RECT  7.755 0.630 7.985 1.385 ;
        RECT  6.455 0.630 6.690 1.170 ;
        RECT  5.300 0.940 6.690 1.170 ;
        RECT  2.120 0.980 2.465 1.415 ;
        RECT  8.810 0.750 9.040 1.385 ;
        RECT  7.755 1.155 9.040 1.385 ;
        RECT  4.085 0.630 4.315 1.410 ;
        RECT  2.120 1.180 4.315 1.410 ;
        RECT  2.120 1.180 2.965 1.415 ;
        RECT  10.140 0.750 10.370 1.500 ;
        RECT  10.340 1.270 10.590 2.145 ;
        RECT  8.520 1.155 8.860 2.085 ;
        RECT  10.340 1.805 10.680 2.145 ;
        RECT  2.735 1.180 2.965 2.670 ;
        RECT  2.075 2.440 2.965 2.670 ;
        RECT  2.075 2.440 2.415 3.625 ;
        RECT  11.110 1.180 11.690 1.410 ;
        RECT  11.345 1.070 11.690 1.410 ;
        RECT  9.720 1.800 10.035 2.845 ;
        RECT  10.975 1.190 11.205 2.845 ;
        RECT  6.950 2.035 7.270 3.005 ;
        RECT  9.720 2.560 11.710 2.845 ;
        RECT  6.950 2.775 9.975 3.005 ;
        RECT  9.270 1.230 9.770 1.570 ;
        RECT  7.050 1.090 7.390 1.805 ;
        RECT  9.260 1.565 9.500 1.685 ;
        RECT  6.490 1.575 7.560 1.805 ;
        RECT  7.415 1.615 8.265 1.845 ;
        RECT  8.035 1.615 8.265 2.545 ;
        RECT  9.260 1.565 9.490 2.545 ;
        RECT  12.110 2.065 13.740 2.405 ;
        RECT  8.035 2.315 9.490 2.545 ;
        RECT  6.490 1.575 6.720 3.465 ;
        RECT  10.215 3.075 12.340 3.305 ;
        RECT  12.110 2.065 12.340 3.305 ;
        RECT  6.490 3.235 10.440 3.465 ;
        RECT  9.385 3.235 10.440 3.490 ;
        RECT  7.045 3.235 7.390 3.585 ;
        RECT  9.385 3.235 9.730 4.030 ;
        RECT  2.755 2.900 3.60 3.130 ;
        RECT  2.120 1.180 3.90 1.410 ;
        RECT  6.950 2.775 8.70 3.005 ;
        RECT  10.215 3.075 11.00 3.305 ;
        RECT  6.490 3.235 9.30 3.465 ;
    END
END MU4IX4

MACRO MU4IX2
    CLASS CORE ;
    FOREIGN MU4IX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.906  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.260 1.165 10.600 1.505 ;
        RECT  10.350 1.165 10.585 3.240 ;
        RECT  10.100 3.260 10.440 4.180 ;
        RECT  10.205 2.860 10.440 4.180 ;
        RECT  10.260 1.165 10.585 1.510 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.676  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.200 1.875 9.955 2.215 ;
        RECT  9.575 1.640 9.955 2.215 ;
        END
    END S1
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.020 2.270 3.665 2.640 ;
        RECT  3.020 2.240 3.380 2.640 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.947  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.250 0.655 2.625 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.505 1.600 6.175 2.035 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.000 1.625 1.340 2.205 ;
        RECT  0.755 1.625 1.340 2.020 ;
        END
    END IN0
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.625 1.640 4.235 2.040 ;
        END
    END IN2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 3.260 11.160 5.280 ;
        RECT  9.380 3.825 9.720 5.280 ;
        RECT  8.215 3.540 8.555 5.280 ;
        RECT  5.810 2.900 6.165 5.280 ;
        RECT  3.320 3.330 3.660 5.280 ;
        RECT  0.935 3.315 1.275 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.820 -0.400 11.160 0.730 ;
        RECT  9.500 -0.400 9.840 0.900 ;
        RECT  8.170 -0.400 8.510 1.405 ;
        RECT  5.785 -0.400 6.130 0.710 ;
        RECT  3.360 -0.400 3.710 0.950 ;
        RECT  0.940 -0.400 1.280 0.915 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.845 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  1.610 1.830 2.175 2.170 ;
        RECT  0.215 2.855 1.840 3.085 ;
        RECT  4.465 1.870 4.695 3.100 ;
        RECT  2.755 2.870 4.695 3.100 ;
        RECT  1.610 1.145 1.840 4.085 ;
        RECT  0.215 2.855 0.555 3.880 ;
        RECT  2.755 2.870 2.985 4.085 ;
        RECT  1.610 3.855 2.985 4.085 ;
        RECT  4.600 1.145 4.990 1.585 ;
        RECT  5.955 2.330 6.240 2.670 ;
        RECT  4.925 2.440 6.240 2.670 ;
        RECT  4.925 1.360 5.155 3.680 ;
        RECT  4.545 3.340 5.155 3.680 ;
        RECT  4.085 0.685 5.515 0.915 ;
        RECT  5.285 0.685 5.515 1.170 ;
        RECT  6.440 0.825 7.845 1.055 ;
        RECT  5.285 0.940 6.675 1.170 ;
        RECT  4.085 0.685 4.315 1.410 ;
        RECT  2.155 1.180 4.315 1.410 ;
        RECT  2.155 1.075 2.500 1.415 ;
        RECT  7.615 0.825 7.845 2.145 ;
        RECT  7.615 1.805 8.315 2.145 ;
        RECT  2.405 1.180 2.635 2.630 ;
        RECT  2.240 2.400 2.470 3.625 ;
        RECT  2.130 2.760 2.470 3.625 ;
        RECT  8.740 1.285 9.270 1.625 ;
        RECT  6.930 2.020 7.220 2.720 ;
        RECT  8.740 1.285 8.970 2.720 ;
        RECT  6.930 2.490 9.315 2.720 ;
        RECT  8.915 2.485 9.315 2.850 ;
        RECT  7.020 1.285 7.360 1.730 ;
        RECT  6.470 1.500 7.360 1.730 ;
        RECT  9.550 2.545 9.975 2.890 ;
        RECT  6.470 1.500 6.700 3.250 ;
        RECT  6.470 2.965 7.400 3.250 ;
        RECT  9.550 2.545 9.780 3.310 ;
        RECT  7.020 3.080 9.780 3.310 ;
        RECT  7.020 2.965 7.365 4.180 ;
        RECT  2.155 1.180 3.20 1.410 ;
        RECT  6.930 2.490 8.70 2.720 ;
        RECT  7.020 3.080 8.70 3.310 ;
    END
END MU4IX2

MACRO MU4IX1
    CLASS CORE ;
    FOREIGN MU4IX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 0.920 10.585 4.180 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.165 1.890 9.955 2.230 ;
        RECT  9.575 1.640 9.955 2.230 ;
        END
    END S1
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.695 2.250 3.480 2.640 ;
        RECT  3.140 1.660 3.480 2.640 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.546  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.205 0.615 2.615 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.600 1.520 6.175 2.020 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.605 1.340 2.020 ;
        END
    END IN0
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.720 1.640 4.290 2.020 ;
        RECT  3.720 1.640 4.060 2.520 ;
        END
    END IN2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 3.575 9.810 5.280 ;
        RECT  8.095 3.540 8.435 5.280 ;
        RECT  5.795 2.960 6.135 5.280 ;
        RECT  3.320 3.480 3.660 5.280 ;
        RECT  0.980 3.305 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.430 -0.400 9.770 0.910 ;
        RECT  8.130 -0.400 8.470 1.540 ;
        RECT  5.745 -0.400 6.090 0.710 ;
        RECT  3.410 -0.400 3.760 0.915 ;
        RECT  0.980 -0.400 1.320 0.915 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.635 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  1.610 1.930 1.955 2.270 ;
        RECT  1.610 1.145 1.840 3.250 ;
        RECT  4.515 2.095 4.855 2.990 ;
        RECT  3.990 2.760 4.855 2.990 ;
        RECT  0.220 2.845 1.840 3.075 ;
        RECT  3.990 2.760 4.220 3.250 ;
        RECT  1.610 3.020 4.220 3.250 ;
        RECT  0.220 2.845 0.580 3.365 ;
        RECT  4.690 1.110 5.030 1.815 ;
        RECT  4.690 1.585 5.315 1.815 ;
        RECT  5.085 2.280 6.280 2.625 ;
        RECT  5.085 1.585 5.315 3.560 ;
        RECT  4.520 3.220 5.315 3.560 ;
        RECT  4.085 0.630 5.515 0.860 ;
        RECT  5.285 0.630 5.515 1.170 ;
        RECT  6.440 0.770 7.845 1.000 ;
        RECT  2.185 0.980 2.550 1.375 ;
        RECT  5.285 0.940 6.675 1.170 ;
        RECT  4.085 0.630 4.315 1.375 ;
        RECT  2.185 1.145 4.315 1.375 ;
        RECT  7.615 0.770 7.845 2.150 ;
        RECT  7.615 1.810 8.230 2.150 ;
        RECT  2.185 0.980 2.465 2.790 ;
        RECT  2.170 2.450 2.465 2.790 ;
        RECT  8.700 1.285 9.270 1.625 ;
        RECT  6.970 1.960 7.310 2.650 ;
        RECT  8.700 1.285 8.930 2.850 ;
        RECT  6.970 2.420 8.930 2.650 ;
        RECT  8.700 2.565 9.195 2.850 ;
        RECT  6.980 1.230 7.320 1.730 ;
        RECT  6.510 1.500 7.320 1.730 ;
        RECT  6.510 1.500 6.740 3.240 ;
        RECT  6.510 2.955 7.285 3.240 ;
        RECT  9.620 2.735 9.960 3.310 ;
        RECT  6.945 3.080 9.960 3.310 ;
        RECT  6.945 2.955 7.285 3.875 ;
        RECT  1.610 3.020 3.60 3.250 ;
        RECT  2.185 1.145 3.50 1.375 ;
        RECT  6.945 3.080 8.80 3.310 ;
    END
END MU4IX1

MACRO MU4IX0
    CLASS CORE ;
    FOREIGN MU4IX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN IN2
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.285 2.530 ;
        END
    END IN2
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.480 2.020 ;
        END
    END IN1
    PIN S0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.405  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.610 0.615 2.030 ;
        END
    END S0
    PIN IN3
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.485 1.640 6.175 1.970 ;
        RECT  5.485 1.640 5.825 2.110 ;
        END
    END IN3
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.255 1.380 2.615 ;
        END
    END IN0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.010 1.640 10.585 2.020 ;
        RECT  10.010 1.170 10.350 3.045 ;
        END
    END Q
    PIN S1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.266  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.290 3.470 8.065 3.850 ;
        END
    END S1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.010 -0.400 10.350 0.710 ;
        RECT  8.280 -0.400 8.625 1.315 ;
        RECT  5.970 -0.400 6.320 0.660 ;
        RECT  3.505 -0.400 3.855 0.915 ;
        RECT  0.980 -0.400 1.320 0.915 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.985 3.505 10.350 5.280 ;
        RECT  8.295 2.965 8.565 5.280 ;
        RECT  8.280 2.965 8.565 3.305 ;
        RECT  5.810 2.850 6.150 5.280 ;
        RECT  3.340 3.285 3.680 5.280 ;
        RECT  1.025 3.305 1.365 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.635 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  1.610 1.930 1.955 2.270 ;
        RECT  1.610 1.145 1.840 3.195 ;
        RECT  2.795 2.760 4.745 2.990 ;
        RECT  4.515 1.555 4.745 2.990 ;
        RECT  0.230 2.845 1.840 3.075 ;
        RECT  1.610 2.965 3.025 3.195 ;
        RECT  0.230 2.845 0.590 3.565 ;
        RECT  4.740 1.090 5.205 1.325 ;
        RECT  6.160 2.250 6.500 2.570 ;
        RECT  4.975 2.340 6.500 2.570 ;
        RECT  4.975 1.090 5.205 3.505 ;
        RECT  4.550 3.220 5.205 3.505 ;
        RECT  4.085 0.630 5.670 0.860 ;
        RECT  6.555 0.630 8.050 0.860 ;
        RECT  5.440 0.630 5.670 1.120 ;
        RECT  6.555 0.630 6.785 1.120 ;
        RECT  5.440 0.890 6.785 1.120 ;
        RECT  2.185 1.000 2.550 1.375 ;
        RECT  4.085 0.630 4.315 1.375 ;
        RECT  2.185 1.145 4.315 1.375 ;
        RECT  7.820 0.630 8.050 1.815 ;
        RECT  7.820 1.545 8.455 1.815 ;
        RECT  2.185 1.000 2.415 2.735 ;
        RECT  2.185 2.450 2.565 2.735 ;
        RECT  7.290 1.855 7.590 2.275 ;
        RECT  9.080 1.010 9.420 2.275 ;
        RECT  7.290 2.045 9.540 2.275 ;
        RECT  9.255 2.045 9.540 2.790 ;
        RECT  7.050 1.090 7.395 1.620 ;
        RECT  6.830 1.390 7.060 2.735 ;
        RECT  6.830 2.505 9.025 2.735 ;
        RECT  8.795 2.505 9.025 3.325 ;
        RECT  7.090 2.505 7.430 3.140 ;
        RECT  8.795 3.020 9.745 3.325 ;
        RECT  2.185 1.145 3.20 1.375 ;
        RECT  7.290 2.045 8.30 2.275 ;
        RECT  6.830 2.505 8.20 2.735 ;
    END
END MU4IX0

MACRO MU2X4
    CLASS CORE ;
    FOREIGN MU2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.877  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.190 2.445 2.390 2.675 ;
        RECT  1.890 2.120 2.390 2.675 ;
        RECT  0.190 2.120 0.530 2.675 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.330  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.770 0.700 6.175 2.025 ;
        RECT  5.780 0.700 6.120 4.180 ;
        RECT  4.450 2.810 6.120 3.040 ;
        RECT  5.770 0.700 6.120 3.040 ;
        RECT  4.450 1.090 6.175 1.425 ;
        RECT  4.340 3.065 4.680 4.180 ;
        RECT  4.450 2.810 4.680 4.180 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.600 2.115 4.285 2.640 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.225 1.690 1.565 2.215 ;
        RECT  0.745 1.690 1.565 2.030 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.020 -0.400 5.360 0.710 ;
        RECT  3.900 -0.400 4.240 0.710 ;
        RECT  0.945 -0.400 1.285 1.000 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.060 3.270 5.400 5.280 ;
        RECT  3.620 3.065 3.965 5.280 ;
        RECT  0.985 3.365 1.325 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.225 0.700 0.565 1.460 ;
        RECT  0.225 1.230 2.295 1.460 ;
        RECT  2.065 1.230 2.295 1.845 ;
        RECT  2.065 1.615 2.910 1.845 ;
        RECT  2.620 1.615 2.910 2.215 ;
        RECT  2.620 1.615 2.850 3.135 ;
        RECT  0.225 2.905 2.850 3.135 ;
        RECT  0.225 2.905 0.565 4.060 ;
        RECT  2.710 1.020 3.370 1.360 ;
        RECT  3.140 1.655 4.765 1.885 ;
        RECT  4.515 1.655 4.765 2.445 ;
        RECT  4.515 2.105 5.540 2.445 ;
        RECT  3.140 1.020 3.370 3.595 ;
        RECT  2.170 3.365 3.370 3.595 ;
        RECT  2.170 3.365 2.510 4.180 ;
        RECT  0.225 1.230 1.50 1.460 ;
        RECT  0.225 2.905 1.10 3.135 ;
    END
END MU2X4

MACRO MU2X2
    CLASS CORE ;
    FOREIGN MU2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.623  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.685 2.405 2.030 2.745 ;
        RECT  1.485 2.480 1.715 3.240 ;
        RECT  0.200 3.710 1.615 3.940 ;
        RECT  1.385 2.860 1.615 3.940 ;
        RECT  0.200 3.710 0.540 4.100 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 1.640 4.915 2.030 ;
        RECT  3.910 2.730 4.745 2.960 ;
        RECT  4.515 1.165 4.745 2.960 ;
        RECT  3.955 1.165 4.745 1.510 ;
        RECT  3.800 3.270 4.140 4.180 ;
        RECT  3.910 2.730 4.140 4.180 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.300 2.220 3.675 2.875 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.720 1.690 1.340 2.215 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.520 -0.400 4.860 0.710 ;
        RECT  3.395 -0.400 3.735 0.710 ;
        RECT  0.980 -0.400 1.320 1.000 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.520 3.270 4.860 5.280 ;
        RECT  3.080 3.250 3.425 5.280 ;
        RECT  0.755 4.185 1.080 5.280 ;
        RECT  0.770 4.170 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.815 0.560 1.460 ;
        RECT  0.180 1.230 1.870 1.460 ;
        RECT  1.640 1.230 1.870 2.130 ;
        RECT  1.640 1.900 2.610 2.130 ;
        RECT  2.325 1.900 2.610 2.280 ;
        RECT  0.180 0.815 0.410 3.480 ;
        RECT  0.180 2.660 0.520 3.480 ;
        RECT  2.205 1.050 3.070 1.390 ;
        RECT  2.840 1.745 4.285 1.975 ;
        RECT  3.945 1.745 4.285 2.240 ;
        RECT  2.840 1.050 3.070 2.775 ;
        RECT  2.360 2.545 3.070 2.775 ;
        RECT  2.360 2.545 2.590 3.300 ;
        RECT  1.945 3.070 2.590 3.300 ;
        RECT  1.945 3.070 2.270 4.045 ;
        RECT  1.930 3.400 2.270 4.045 ;
    END
END MU2X2

MACRO MU2X1
    CLASS CORE ;
    FOREIGN MU2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.347  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.165 1.145 2.680 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.185 2.860 4.915 3.240 ;
        RECT  4.510 1.160 4.740 3.240 ;
        RECT  4.185 2.860 4.525 3.770 ;
        RECT  4.390 1.160 4.740 1.505 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 2.205 3.760 2.670 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 1.690 1.770 2.215 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.670 -0.400 4.010 1.465 ;
        RECT  1.170 -0.400 1.510 1.000 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.455 2.900 3.800 5.280 ;
        RECT  1.100 2.940 1.440 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.285 1.130 0.710 1.460 ;
        RECT  0.285 1.230 2.230 1.460 ;
        RECT  2.000 1.230 2.230 2.240 ;
        RECT  2.000 1.900 2.505 2.240 ;
        RECT  0.285 1.130 0.520 3.255 ;
        RECT  0.285 2.915 0.720 3.255 ;
        RECT  2.460 1.145 3.075 1.485 ;
        RECT  2.845 1.745 4.280 1.975 ;
        RECT  3.990 1.745 4.280 2.240 ;
        RECT  2.845 1.145 3.075 3.250 ;
        RECT  2.250 3.020 3.075 3.250 ;
        RECT  2.250 3.020 2.590 3.370 ;
    END
END MU2X1

MACRO MU2X0
    CLASS CORE ;
    FOREIGN MU2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.266  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.610 0.625 1.995 ;
        RECT  0.120 1.610 0.565 2.115 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.449  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.825 2.860 4.285 3.250 ;
        RECT  3.940 1.360 4.285 3.250 ;
        RECT  3.890 1.360 4.285 1.700 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.640 3.655 2.020 ;
        RECT  2.780 1.470 3.110 2.020 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.139  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.245 1.330 2.650 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.290 -0.400 3.645 1.060 ;
        RECT  0.980 -0.400 1.320 0.915 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.200 3.510 3.540 5.280 ;
        RECT  0.980 3.340 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.635 0.520 1.375 ;
        RECT  0.180 1.145 1.840 1.375 ;
        RECT  1.610 2.225 1.995 2.565 ;
        RECT  1.610 1.145 1.840 3.110 ;
        RECT  0.180 2.880 1.840 3.110 ;
        RECT  0.180 2.880 0.520 3.620 ;
        RECT  2.210 1.280 2.550 1.620 ;
        RECT  2.225 1.280 2.550 2.620 ;
        RECT  2.225 2.280 3.710 2.620 ;
        RECT  2.225 1.280 2.510 4.000 ;
        RECT  2.170 3.660 2.510 4.000 ;
    END
END MU2X0

MACRO MU2IX4
    CLASS CORE ;
    FOREIGN MU2IX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 1.083  LAYER MET1  ;
        ANTENNAGATEAREA 2.034  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.815 3.710 13.375 4.050 ;
        RECT  12.815 2.450 13.045 4.050 ;
        RECT  11.090 2.450 13.045 2.680 ;
        RECT  11.090 2.340 11.375 2.680 ;
        RECT  2.435 2.340 2.720 2.710 ;
        RECT  1.625 2.480 2.720 2.710 ;
        RECT  0.750 2.540 1.800 2.770 ;
        RECT  0.750 2.540 0.980 3.700 ;
        RECT  0.125 3.470 0.760 4.050 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.701  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.305 1.145 12.645 1.670 ;
        RECT  9.155 1.145 12.645 1.375 ;
        RECT  10.300 3.370 11.395 3.600 ;
        RECT  3.370 3.305 10.465 3.535 ;
        RECT  9.155 1.035 9.715 1.375 ;
        RECT  4.420 1.515 9.385 1.745 ;
        RECT  9.155 1.035 9.385 1.745 ;
        RECT  6.905 0.880 7.245 1.745 ;
        RECT  3.905 3.250 5.780 3.535 ;
        RECT  5.550 1.515 5.780 3.535 ;
        RECT  4.420 1.040 4.650 1.745 ;
        RECT  1.135 1.150 4.650 1.380 ;
        RECT  4.090 1.040 4.650 1.380 ;
        RECT  3.905 2.860 4.285 3.535 ;
        RECT  2.425 3.400 3.560 3.585 ;
        RECT  2.425 3.400 3.515 3.630 ;
        RECT  1.135 1.150 1.475 1.790 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.584  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.660 1.975 7.560 2.615 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.584  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.970 3.830 11.855 4.060 ;
        RECT  11.625 2.910 11.855 4.060 ;
        RECT  10.630 2.910 11.855 3.140 ;
        RECT  10.630 2.065 10.860 3.140 ;
        RECT  10.205 2.065 10.860 2.630 ;
        RECT  3.705 3.765 10.135 3.995 ;
        RECT  1.965 3.860 3.895 4.090 ;
        RECT  2.950 2.070 3.520 2.355 ;
        RECT  1.965 2.940 3.180 3.170 ;
        RECT  2.950 2.070 3.180 3.170 ;
        RECT  1.965 2.940 2.195 4.090 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.035 -0.400 13.375 0.710 ;
        RECT  10.565 -0.400 11.455 0.915 ;
        RECT  8.225 -0.400 8.565 1.285 ;
        RECT  5.585 -0.400 5.925 1.285 ;
        RECT  2.365 -0.400 3.240 0.920 ;
        RECT  0.485 -0.400 0.825 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.245 2.910 12.585 5.280 ;
        RECT  9.465 4.225 9.805 5.280 ;
        RECT  6.940 4.225 7.280 5.280 ;
        RECT  4.085 4.225 4.425 5.280 ;
        RECT  1.235 3.000 1.575 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.745 1.610 4.190 1.840 ;
        RECT  0.445 1.090 0.785 2.310 ;
        RECT  0.445 2.020 1.975 2.250 ;
        RECT  1.745 1.610 1.975 2.250 ;
        RECT  0.180 2.080 1.390 2.310 ;
        RECT  3.850 1.610 4.190 2.570 ;
        RECT  3.850 2.340 5.320 2.570 ;
        RECT  5.035 2.340 5.320 2.680 ;
        RECT  0.180 2.080 0.520 3.240 ;
        RECT  9.615 1.605 12.075 1.835 ;
        RECT  11.845 1.605 12.075 2.130 ;
        RECT  11.845 1.900 13.615 2.130 ;
        RECT  13.075 1.090 13.415 2.220 ;
        RECT  12.310 1.900 13.615 2.220 ;
        RECT  9.615 1.605 9.955 2.680 ;
        RECT  8.110 2.340 9.955 2.680 ;
        RECT  6.010 2.340 6.295 3.075 ;
        RECT  8.110 2.340 8.340 3.075 ;
        RECT  6.010 2.845 8.340 3.075 ;
        RECT  13.275 1.900 13.615 3.240 ;
        RECT  1.745 1.610 3.40 1.840 ;
        RECT  9.615 1.605 11.80 1.835 ;
        RECT  6.010 2.845 7.40 3.075 ;
    END
END MU2IX4

MACRO MU2IX2
    CLASS CORE ;
    FOREIGN MU2IX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.704  LAYER MET1  ;
        ANTENNAGATEAREA 1.091  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.575 3.460 7.140 3.800 ;
        RECT  6.575 2.450 6.805 3.800 ;
        RECT  5.560 2.450 6.805 2.680 ;
        RECT  5.560 2.340 5.875 2.680 ;
        RECT  0.900 2.450 1.975 2.680 ;
        RECT  1.685 2.340 1.975 2.680 ;
        RECT  0.900 2.450 1.135 3.240 ;
        RECT  0.420 3.475 0.985 3.800 ;
        RECT  0.755 2.860 0.985 3.800 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.330  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.640 3.450 5.140 3.790 ;
        RECT  4.155 0.850 5.140 1.190 ;
        RECT  4.640 3.010 4.870 3.790 ;
        RECT  2.690 3.010 4.870 3.240 ;
        RECT  3.905 2.860 4.385 3.240 ;
        RECT  4.155 0.850 4.385 3.240 ;
        RECT  3.150 1.750 4.385 1.980 ;
        RECT  3.150 0.850 3.380 1.980 ;
        RECT  2.420 0.850 3.380 1.190 ;
        RECT  2.420 3.450 2.920 3.790 ;
        RECT  2.690 3.010 2.920 3.790 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.925 2.630 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.220 1.880 6.560 2.220 ;
        RECT  5.100 1.880 6.560 2.110 ;
        RECT  5.395 3.470 6.175 3.850 ;
        RECT  4.180 4.020 5.625 4.250 ;
        RECT  5.395 2.910 5.625 4.250 ;
        RECT  5.100 2.910 5.625 3.140 ;
        RECT  5.100 1.880 5.330 3.140 ;
        RECT  4.180 3.470 4.410 4.250 ;
        RECT  3.150 3.470 4.410 3.700 ;
        RECT  1.960 4.020 3.380 4.250 ;
        RECT  3.150 3.470 3.380 4.250 ;
        RECT  1.960 2.910 2.435 3.140 ;
        RECT  2.205 1.880 2.435 3.140 ;
        RECT  1.000 1.880 2.435 2.110 ;
        RECT  1.960 2.910 2.190 4.250 ;
        RECT  1.000 1.880 1.340 2.220 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.240 -0.400 6.580 1.165 ;
        RECT  3.610 -0.400 3.925 1.520 ;
        RECT  0.980 -0.400 1.320 1.165 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.480 4.065 6.820 5.280 ;
        RECT  3.610 3.930 3.950 5.280 ;
        RECT  0.740 4.065 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.825 0.520 1.650 ;
        RECT  0.180 1.420 2.895 1.650 ;
        RECT  2.665 1.420 2.895 2.680 ;
        RECT  2.665 2.340 3.000 2.680 ;
        RECT  0.180 0.825 0.410 3.245 ;
        RECT  0.180 2.915 0.520 3.245 ;
        RECT  4.615 1.420 7.380 1.650 ;
        RECT  4.615 1.420 4.870 2.680 ;
        RECT  7.040 0.825 7.380 3.230 ;
        RECT  0.180 1.420 1.40 1.650 ;
        RECT  4.615 1.420 6.30 1.650 ;
    END
END MU2IX2

MACRO MU2IX1
    CLASS CORE ;
    FOREIGN MU2IX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.551  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.575 2.340 2.030 2.675 ;
        RECT  1.575 2.340 1.810 3.240 ;
        RECT  0.420 3.475 1.615 3.800 ;
        RECT  1.385 2.860 1.615 3.800 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.364  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.865 1.415 3.095 2.665 ;
        RECT  2.260 2.520 3.065 2.750 ;
        RECT  2.795 1.030 3.025 1.650 ;
        RECT  2.110 1.030 3.025 1.410 ;
        RECT  2.260 2.520 2.490 3.135 ;
        RECT  2.040 2.905 2.380 4.180 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 2.035 3.665 2.705 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.392  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.050 1.340 2.390 ;
        RECT  0.755 2.050 1.135 2.630 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.260 -0.400 3.600 1.250 ;
        RECT  0.960 -0.400 1.300 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.190 2.955 3.530 5.280 ;
        RECT  0.740 4.030 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.590 1.800 1.820 ;
        RECT  1.570 1.590 1.800 2.110 ;
        RECT  1.570 1.880 2.635 2.110 ;
        RECT  2.350 1.880 2.635 2.290 ;
        RECT  0.180 1.140 0.520 3.245 ;
    END
END MU2IX1

MACRO MU2IX0
    CLASS CORE ;
    FOREIGN MU2IX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.276  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.640 0.625 2.010 ;
        RECT  0.120 1.640 0.565 2.125 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.726  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.170 2.860 2.550 3.675 ;
        RECT  2.185 1.000 2.550 3.675 ;
        RECT  2.015 2.860 2.550 3.250 ;
        END
    END Q
    PIN IN1
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.115 2.185 3.655 2.630 ;
        END
    END IN1
    PIN IN0
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.255 1.320 2.640 ;
        END
    END IN0
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.260 -0.400 3.615 0.760 ;
        RECT  0.980 -0.400 1.320 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.210 3.650 3.550 5.280 ;
        RECT  1.015 3.335 1.355 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.635 0.520 1.410 ;
        RECT  0.180 1.180 1.780 1.410 ;
        RECT  1.550 1.850 1.955 2.215 ;
        RECT  1.550 1.180 1.780 3.105 ;
        RECT  0.215 2.875 1.780 3.105 ;
        RECT  0.215 2.875 0.555 3.675 ;
    END
END MU2IX0

MACRO LSOGCPX8
    CLASS CORE ;
    FOREIGN LSOGCPX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.380 1.105 18.775 3.740 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.800 11.845 2.630 ;
        RECT  10.935 1.800 11.845 2.140 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.795 2.060 16.275 2.630 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.142  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.155 2.660 3.505 4.180 ;
        RECT  3.155 0.725 3.505 1.700 ;
        RECT  3.155 0.725 3.435 4.180 ;
        RECT  0.125 2.090 3.435 2.430 ;
        RECT  1.725 2.090 2.070 4.180 ;
        RECT  1.725 0.725 2.065 4.180 ;
        RECT  0.125 0.725 0.625 4.180 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.444  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.150 1.640 8.695 2.430 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  17.660 2.820 18.000 5.280 ;
        RECT  16.175 3.315 16.515 5.280 ;
        RECT  12.855 3.565 14.215 5.280 ;
        RECT  11.820 3.705 12.160 5.280 ;
        RECT  9.690 3.580 10.030 5.280 ;
        RECT  8.205 3.120 8.545 5.280 ;
        RECT  6.765 2.760 7.105 5.280 ;
        RECT  5.325 2.760 5.665 5.280 ;
        RECT  3.885 2.760 4.225 5.280 ;
        RECT  2.445 2.660 2.785 5.280 ;
        RECT  1.005 2.660 1.345 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  17.660 -0.400 18.000 1.495 ;
        RECT  16.160 -0.400 16.500 1.025 ;
        RECT  13.980 -0.400 14.320 1.670 ;
        RECT  11.780 -0.400 12.120 0.970 ;
        RECT  10.360 -0.400 10.700 0.970 ;
        RECT  9.050 -0.400 9.390 1.560 ;
        RECT  6.760 -0.400 7.100 1.490 ;
        RECT  3.885 -0.400 4.760 1.700 ;
        RECT  2.445 -0.400 2.785 1.705 ;
        RECT  1.005 -0.400 1.345 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  7.485 1.090 8.250 1.410 ;
        RECT  5.610 1.125 5.950 2.270 ;
        RECT  3.695 1.930 7.825 2.270 ;
        RECT  7.485 2.660 9.265 2.890 ;
        RECT  4.605 1.930 4.945 3.680 ;
        RECT  6.045 1.930 6.390 3.680 ;
        RECT  7.485 1.090 7.825 3.680 ;
        RECT  8.925 2.660 9.265 3.680 ;
        RECT  9.620 1.350 10.100 1.690 ;
        RECT  9.170 1.900 9.850 2.240 ;
        RECT  9.620 1.350 9.850 3.115 ;
        RECT  9.620 2.830 10.590 3.115 ;
        RECT  10.475 1.280 11.500 1.570 ;
        RECT  10.110 1.950 10.705 2.290 ;
        RECT  10.475 1.280 10.705 2.600 ;
        RECT  10.475 2.370 11.050 2.600 ;
        RECT  10.820 2.370 11.050 4.010 ;
        RECT  10.670 3.650 11.050 4.010 ;
        RECT  12.580 0.630 12.920 2.215 ;
        RECT  12.580 1.875 13.290 2.215 ;
        RECT  12.580 0.630 12.830 3.335 ;
        RECT  14.550 2.740 15.105 3.080 ;
        RECT  12.110 2.765 12.830 3.105 ;
        RECT  14.550 2.740 14.780 3.335 ;
        RECT  12.575 3.105 14.780 3.335 ;
        RECT  13.180 1.305 13.750 1.645 ;
        RECT  13.520 1.305 13.750 2.875 ;
        RECT  13.520 2.070 15.105 2.410 ;
        RECT  13.520 2.070 13.770 2.875 ;
        RECT  13.430 2.590 13.770 2.875 ;
        RECT  15.170 1.420 16.730 1.760 ;
        RECT  15.335 1.420 16.730 1.770 ;
        RECT  15.335 1.420 15.565 3.695 ;
        RECT  15.025 3.355 15.565 3.695 ;
        RECT  16.960 0.910 17.300 4.250 ;
        RECT  16.960 3.905 17.425 4.250 ;
        RECT  3.695 1.930 6.20 2.270 ;
        RECT  12.575 3.105 13.50 3.335 ;
    END
END LSOGCPX8

MACRO LSOGCPX6
    CLASS CORE ;
    FOREIGN LSOGCPX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 1.105 16.885 3.740 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 1.800 9.955 2.630 ;
        RECT  9.045 1.800 9.955 2.140 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.905 2.060 14.390 2.630 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.689  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 0.790 2.680 4.180 ;
        RECT  0.900 2.090 2.680 2.430 ;
        RECT  0.900 2.090 1.245 4.180 ;
        RECT  0.900 0.790 1.240 4.180 ;
        RECT  0.755 2.250 1.245 2.630 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.120  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.260 1.640 6.805 2.430 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 2.820 16.110 5.280 ;
        RECT  14.285 3.315 14.625 5.280 ;
        RECT  10.965 3.565 12.325 5.280 ;
        RECT  9.930 3.705 10.270 5.280 ;
        RECT  7.800 3.580 8.140 5.280 ;
        RECT  6.315 3.120 6.655 5.280 ;
        RECT  4.875 2.760 5.215 5.280 ;
        RECT  3.250 2.760 3.590 5.280 ;
        RECT  1.620 2.760 1.960 5.280 ;
        RECT  0.180 2.760 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.770 -0.400 16.110 1.495 ;
        RECT  14.270 -0.400 14.610 1.025 ;
        RECT  12.090 -0.400 12.430 1.670 ;
        RECT  9.890 -0.400 10.230 0.970 ;
        RECT  8.470 -0.400 8.810 0.970 ;
        RECT  7.170 -0.400 7.500 1.520 ;
        RECT  4.870 -0.400 5.210 1.490 ;
        RECT  3.060 -0.400 3.400 1.130 ;
        RECT  1.620 -0.400 1.960 1.705 ;
        RECT  0.180 -0.400 0.520 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  5.595 1.090 6.360 1.410 ;
        RECT  3.720 1.380 4.060 2.270 ;
        RECT  2.940 1.930 5.935 2.270 ;
        RECT  5.595 2.660 7.375 2.890 ;
        RECT  4.155 1.930 4.500 3.680 ;
        RECT  5.595 1.090 5.935 3.680 ;
        RECT  7.035 2.660 7.375 3.680 ;
        RECT  7.730 1.350 8.210 1.690 ;
        RECT  7.280 1.900 7.960 2.240 ;
        RECT  7.730 1.350 7.960 3.115 ;
        RECT  7.730 2.830 8.700 3.115 ;
        RECT  8.585 1.280 9.610 1.570 ;
        RECT  8.220 1.950 8.815 2.290 ;
        RECT  8.585 1.280 8.815 2.600 ;
        RECT  8.585 2.370 9.160 2.600 ;
        RECT  8.930 2.370 9.160 4.010 ;
        RECT  8.780 3.650 9.160 4.010 ;
        RECT  10.645 0.630 11.030 2.215 ;
        RECT  10.645 1.875 11.400 2.215 ;
        RECT  10.645 0.630 10.875 3.335 ;
        RECT  12.660 2.740 13.215 3.080 ;
        RECT  10.220 2.765 10.875 3.105 ;
        RECT  12.660 2.740 12.890 3.335 ;
        RECT  10.645 3.105 12.890 3.335 ;
        RECT  11.290 1.305 11.860 1.645 ;
        RECT  11.630 1.305 11.860 2.875 ;
        RECT  11.630 2.070 13.215 2.410 ;
        RECT  11.630 2.070 11.880 2.875 ;
        RECT  11.540 2.590 11.880 2.875 ;
        RECT  13.280 1.420 14.840 1.760 ;
        RECT  13.445 1.420 14.840 1.770 ;
        RECT  13.445 1.420 13.675 3.695 ;
        RECT  13.135 3.355 13.675 3.695 ;
        RECT  15.070 0.910 15.410 4.250 ;
        RECT  15.070 3.900 15.535 4.250 ;
        RECT  2.940 1.930 4.00 2.270 ;
        RECT  10.645 3.105 11.40 3.335 ;
    END
END LSOGCPX6

MACRO LSOGCPX4
    CLASS CORE ;
    FOREIGN LSOGCPX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 1.105 14.365 3.740 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.800 7.435 2.630 ;
        RECT  6.525 1.800 7.435 2.140 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.385 2.060 11.865 2.630 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.254  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 2.760 1.975 4.010 ;
        RECT  1.620 1.145 1.970 1.485 ;
        RECT  1.620 1.145 1.930 4.010 ;
        RECT  1.385 2.220 1.930 2.630 ;
        RECT  0.190 2.220 1.930 2.530 ;
        RECT  0.190 1.140 0.560 2.530 ;
        RECT  0.190 1.140 0.535 4.010 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.796  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.740 1.640 4.285 2.430 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.250 2.820 13.590 5.280 ;
        RECT  11.765 3.315 12.105 5.280 ;
        RECT  8.445 3.565 9.805 5.280 ;
        RECT  7.410 3.705 7.750 5.280 ;
        RECT  5.280 3.580 5.620 5.280 ;
        RECT  3.795 3.120 4.135 5.280 ;
        RECT  2.355 2.760 2.695 5.280 ;
        RECT  0.915 2.835 1.255 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.250 -0.400 13.590 1.495 ;
        RECT  11.750 -0.400 12.090 1.025 ;
        RECT  9.570 -0.400 9.910 1.670 ;
        RECT  7.370 -0.400 7.710 0.970 ;
        RECT  5.950 -0.400 6.290 0.970 ;
        RECT  4.640 -0.400 4.980 1.560 ;
        RECT  2.350 -0.400 2.690 1.490 ;
        RECT  0.910 -0.400 1.260 1.485 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.075 1.090 3.840 1.410 ;
        RECT  2.160 2.135 3.415 2.475 ;
        RECT  3.075 2.660 4.855 2.890 ;
        RECT  3.075 1.090 3.415 3.680 ;
        RECT  4.515 2.660 4.855 3.680 ;
        RECT  5.210 1.350 5.690 1.690 ;
        RECT  4.760 1.900 5.440 2.240 ;
        RECT  5.210 1.350 5.440 3.115 ;
        RECT  5.210 2.830 6.180 3.115 ;
        RECT  6.065 1.280 7.090 1.570 ;
        RECT  5.700 1.950 6.295 2.290 ;
        RECT  6.065 1.280 6.295 2.600 ;
        RECT  6.065 2.370 6.640 2.600 ;
        RECT  6.410 2.370 6.640 4.010 ;
        RECT  6.260 3.650 6.640 4.010 ;
        RECT  8.170 1.875 8.790 2.215 ;
        RECT  8.170 0.630 8.510 3.335 ;
        RECT  10.140 2.740 10.695 3.080 ;
        RECT  7.700 2.780 8.510 3.120 ;
        RECT  10.140 2.740 10.370 3.335 ;
        RECT  8.125 3.105 10.370 3.335 ;
        RECT  8.770 1.305 9.340 1.645 ;
        RECT  9.020 1.305 9.340 2.875 ;
        RECT  9.020 2.070 10.695 2.410 ;
        RECT  9.020 2.070 9.360 2.875 ;
        RECT  10.760 1.420 12.320 1.760 ;
        RECT  10.925 1.420 12.320 1.765 ;
        RECT  10.925 1.420 11.155 3.695 ;
        RECT  10.615 3.355 11.155 3.695 ;
        RECT  12.550 0.910 12.890 4.250 ;
        RECT  12.550 3.910 13.015 4.250 ;
        RECT  8.125 3.105 9.80 3.335 ;
    END
END LSOGCPX4

MACRO LSOGCPX3
    CLASS CORE ;
    FOREIGN LSOGCPX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 1.105 12.475 3.740 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.635 2.250 5.545 2.630 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.495 2.060 9.975 2.630 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.345  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.760 1.240 4.180 ;
        RECT  0.755 0.790 1.240 1.700 ;
        RECT  0.755 0.790 1.020 4.180 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.634  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.075 2.285 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.360 2.820 11.700 5.280 ;
        RECT  9.875 3.315 10.215 5.280 ;
        RECT  6.555 3.565 7.915 5.280 ;
        RECT  5.270 3.705 5.610 5.280 ;
        RECT  3.060 3.715 3.400 5.280 ;
        RECT  1.620 3.435 1.960 5.280 ;
        RECT  0.180 2.760 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.360 -0.400 11.700 1.495 ;
        RECT  9.860 -0.400 10.200 1.025 ;
        RECT  7.680 -0.400 8.020 1.670 ;
        RECT  5.380 -0.400 5.720 0.970 ;
        RECT  3.960 -0.400 4.300 0.970 ;
        RECT  1.620 -0.400 1.960 1.080 ;
        RECT  0.180 -0.400 0.520 1.705 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.770 0.700 3.110 1.040 ;
        RECT  2.170 1.180 3.075 1.410 ;
        RECT  2.770 0.700 3.075 1.410 ;
        RECT  1.490 1.310 2.380 1.540 ;
        RECT  1.250 2.185 1.720 2.525 ;
        RECT  1.490 1.310 1.720 3.205 ;
        RECT  1.490 2.975 2.680 3.205 ;
        RECT  2.340 2.975 2.680 4.180 ;
        RECT  3.310 1.370 3.700 1.710 ;
        RECT  1.950 2.240 2.260 2.745 ;
        RECT  3.310 1.370 3.540 2.750 ;
        RECT  1.950 2.515 3.540 2.745 ;
        RECT  3.310 2.520 3.945 2.750 ;
        RECT  3.660 2.520 3.945 3.100 ;
        RECT  4.175 1.280 5.100 1.620 ;
        RECT  3.810 1.950 4.405 2.290 ;
        RECT  4.175 1.280 4.405 4.010 ;
        RECT  4.065 3.650 4.405 4.010 ;
        RECT  6.180 1.275 6.520 2.215 ;
        RECT  6.180 1.875 6.990 2.215 ;
        RECT  6.180 1.275 6.465 3.335 ;
        RECT  8.250 2.740 8.805 3.080 ;
        RECT  5.810 2.765 6.465 3.105 ;
        RECT  8.250 2.740 8.480 3.335 ;
        RECT  6.180 3.105 8.480 3.335 ;
        RECT  6.880 1.305 7.450 1.645 ;
        RECT  7.220 1.305 7.450 2.875 ;
        RECT  7.220 2.070 8.805 2.410 ;
        RECT  7.220 2.070 7.470 2.875 ;
        RECT  7.130 2.590 7.470 2.875 ;
        RECT  8.870 1.420 10.430 1.760 ;
        RECT  9.035 1.420 10.430 1.770 ;
        RECT  9.035 1.420 9.265 3.695 ;
        RECT  8.725 3.355 9.265 3.695 ;
        RECT  10.660 0.910 11.000 4.250 ;
        RECT  10.660 3.910 11.125 4.250 ;
        RECT  6.180 3.105 7.40 3.335 ;
    END
END LSOGCPX3

MACRO LSOGCPX2
    CLASS CORE ;
    FOREIGN LSOGCPX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 1.105 12.475 3.740 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.985 3.445 5.570 3.875 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.495 2.030 9.975 2.630 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.810 1.240 3.240 ;
        RECT  0.850 1.230 1.240 1.570 ;
        RECT  0.850 1.230 1.080 3.240 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 1.630 3.080 2.175 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.360 2.820 11.700 5.280 ;
        RECT  9.875 3.315 10.215 5.280 ;
        RECT  6.555 3.565 7.915 5.280 ;
        RECT  3.425 3.455 4.420 5.280 ;
        RECT  1.515 3.070 1.960 3.425 ;
        RECT  1.515 3.070 1.805 5.280 ;
        RECT  0.150 2.810 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.360 -0.400 11.700 1.495 ;
        RECT  9.860 -0.400 10.200 1.025 ;
        RECT  7.680 -0.400 8.020 1.670 ;
        RECT  5.380 -0.400 5.720 0.970 ;
        RECT  3.960 -0.400 4.300 0.970 ;
        RECT  1.460 -0.400 1.800 0.710 ;
        RECT  0.180 -0.400 0.520 1.575 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.640 0.940 2.990 1.280 ;
        RECT  1.640 0.940 1.870 2.750 ;
        RECT  1.310 2.235 1.870 2.575 ;
        RECT  1.640 2.520 2.420 2.750 ;
        RECT  2.190 2.520 2.420 3.600 ;
        RECT  2.190 3.260 2.680 3.600 ;
        RECT  3.310 1.305 3.700 1.645 ;
        RECT  3.310 1.305 3.580 2.925 ;
        RECT  3.310 2.585 3.860 2.925 ;
        RECT  2.910 2.695 3.860 2.925 ;
        RECT  2.910 2.695 3.195 4.135 ;
        RECT  2.035 3.905 3.195 4.135 ;
        RECT  2.035 3.905 2.320 4.250 ;
        RECT  4.350 1.280 5.100 1.620 ;
        RECT  3.810 1.950 4.580 2.290 ;
        RECT  4.350 1.280 4.580 2.925 ;
        RECT  4.350 2.585 5.610 2.925 ;
        RECT  6.180 1.945 6.900 2.285 ;
        RECT  8.250 2.740 8.805 3.080 ;
        RECT  6.180 1.275 6.520 3.335 ;
        RECT  8.250 2.740 8.480 3.335 ;
        RECT  5.810 3.105 8.480 3.335 ;
        RECT  5.810 3.105 6.150 3.640 ;
        RECT  6.880 1.305 7.450 1.645 ;
        RECT  7.130 1.305 7.450 2.875 ;
        RECT  7.130 2.070 8.805 2.410 ;
        RECT  7.130 2.070 7.470 2.875 ;
        RECT  8.870 1.420 10.430 1.760 ;
        RECT  9.035 1.420 10.430 1.770 ;
        RECT  9.035 1.420 9.265 3.695 ;
        RECT  8.725 3.355 9.265 3.695 ;
        RECT  10.660 0.910 11.000 4.250 ;
        RECT  10.660 3.905 11.125 4.250 ;
        RECT  5.810 3.105 7.90 3.335 ;
    END
END LSOGCPX2

MACRO LSOGCPX1
    CLASS CORE ;
    FOREIGN LSOGCPX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.520 3.560 ;
        RECT  0.125 1.030 0.520 1.370 ;
        RECT  0.125 1.030 0.355 3.560 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.310  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.640 2.030 2.020 ;
        END
    END CLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.510 2.250 9.325 2.630 ;
        RECT  8.510 1.940 8.845 2.630 ;
        END
    END E
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.820 1.360 11.215 3.740 ;
        RECT  10.465 1.360 11.215 1.700 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.845 3.410 4.345 3.910 ;
        END
    END SE
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.260 4.140 10.600 5.280 ;
        RECT  8.905 3.650 9.245 5.280 ;
        RECT  5.455 3.565 6.905 5.280 ;
        RECT  2.705 3.455 3.045 5.280 ;
        RECT  0.820 2.980 1.240 3.335 ;
        RECT  0.820 2.980 1.125 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.465 -0.400 10.805 0.980 ;
        RECT  8.745 -0.400 9.085 1.040 ;
        RECT  6.580 -0.400 6.905 1.670 ;
        RECT  4.490 -0.400 4.830 0.970 ;
        RECT  3.070 -0.400 3.410 0.970 ;
        RECT  0.940 -0.400 1.280 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.510 0.630 2.310 0.980 ;
        RECT  0.750 0.940 1.740 1.170 ;
        RECT  0.590 1.695 0.980 2.030 ;
        RECT  0.750 0.940 0.980 2.750 ;
        RECT  0.750 2.520 1.700 2.750 ;
        RECT  1.470 2.520 1.700 3.335 ;
        RECT  1.470 2.995 1.960 3.335 ;
        RECT  2.370 1.305 2.810 1.645 ;
        RECT  2.370 1.305 2.600 2.925 ;
        RECT  2.370 2.585 2.760 2.925 ;
        RECT  2.190 2.695 2.475 4.035 ;
        RECT  1.355 3.690 2.475 4.035 ;
        RECT  2.830 1.950 4.210 2.290 ;
        RECT  3.870 1.280 4.210 2.925 ;
        RECT  3.870 2.585 4.510 2.925 ;
        RECT  5.765 1.305 6.350 1.645 ;
        RECT  6.030 1.305 6.350 2.875 ;
        RECT  6.030 2.070 7.815 2.410 ;
        RECT  6.030 2.070 6.370 2.875 ;
        RECT  5.290 0.630 5.630 0.950 ;
        RECT  5.290 1.945 5.800 2.285 ;
        RECT  7.240 2.740 7.820 3.080 ;
        RECT  5.290 0.630 5.520 3.335 ;
        RECT  7.240 2.740 7.470 3.335 ;
        RECT  4.710 3.105 7.470 3.335 ;
        RECT  4.710 3.105 5.050 3.640 ;
        RECT  7.755 1.270 9.305 1.610 ;
        RECT  7.755 1.270 8.280 1.760 ;
        RECT  8.050 1.270 8.280 3.695 ;
        RECT  7.715 3.355 8.280 3.695 ;
        RECT  9.555 0.700 9.885 4.145 ;
        RECT  9.475 2.830 9.885 4.145 ;
        RECT  4.710 3.105 6.40 3.335 ;
    END
END LSOGCPX1

MACRO LSOGCPX0
    CLASS CORE ;
    FOREIGN LSOGCPX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.540 2.400 2.180 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.300 0.520 2.980 ;
        RECT  0.125 1.150 0.520 1.490 ;
        RECT  0.125 2.265 0.500 2.980 ;
        RECT  0.125 1.150 0.355 2.980 ;
        END
    END GCLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.665 2.250 9.325 2.630 ;
        RECT  8.665 1.715 8.990 2.630 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.445 1.880 5.020 2.220 ;
        RECT  4.570 1.675 5.020 2.220 ;
        RECT  4.535 1.690 5.020 2.220 ;
        END
    END SE
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.705 2.250 11.215 2.980 ;
        RECT  10.705 1.170 11.155 2.980 ;
        END
    END CGOBS
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.705 3.440 11.045 5.280 ;
        RECT  8.980 3.510 9.320 5.280 ;
        RECT  5.635 3.565 6.905 5.280 ;
        RECT  3.095 3.285 3.435 5.280 ;
        RECT  0.980 2.640 1.320 2.980 ;
        RECT  0.980 2.640 1.285 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.815 -0.400 11.155 0.710 ;
        RECT  9.130 -0.400 9.510 1.025 ;
        RECT  7.005 -0.400 7.435 0.970 ;
        RECT  4.705 -0.400 5.125 0.970 ;
        RECT  3.380 -0.400 3.720 0.970 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.555 0.630 2.350 0.970 ;
        RECT  0.630 1.735 1.785 2.075 ;
        RECT  1.555 0.630 1.785 3.060 ;
        RECT  1.555 2.775 2.120 3.060 ;
        RECT  2.635 1.305 2.920 1.645 ;
        RECT  2.580 2.585 2.920 2.925 ;
        RECT  2.580 2.585 2.865 3.520 ;
        RECT  2.635 1.305 2.865 3.520 ;
        RECT  1.515 3.290 2.865 3.520 ;
        RECT  1.515 3.290 1.800 3.635 ;
        RECT  3.970 1.180 4.390 1.480 ;
        RECT  3.095 2.065 3.380 2.405 ;
        RECT  3.095 2.175 4.200 2.405 ;
        RECT  3.970 1.180 4.200 2.920 ;
        RECT  3.970 2.585 4.760 2.870 ;
        RECT  3.970 2.585 4.750 2.920 ;
        RECT  5.550 1.215 5.865 1.555 ;
        RECT  5.585 1.215 5.865 3.335 ;
        RECT  5.585 1.945 6.110 2.285 ;
        RECT  5.585 1.945 5.870 3.335 ;
        RECT  7.490 2.820 7.860 3.105 ;
        RECT  4.890 3.105 7.850 3.135 ;
        RECT  4.890 3.105 7.720 3.335 ;
        RECT  4.890 3.105 5.175 3.710 ;
        RECT  4.835 3.370 5.175 3.710 ;
        RECT  6.205 1.215 6.625 1.555 ;
        RECT  6.340 1.215 6.625 2.875 ;
        RECT  7.670 2.150 7.955 2.490 ;
        RECT  6.340 2.260 7.955 2.490 ;
        RECT  6.340 2.260 6.630 2.875 ;
        RECT  6.290 2.590 6.630 2.875 ;
        RECT  8.090 1.255 9.515 1.485 ;
        RECT  8.090 1.255 8.415 1.650 ;
        RECT  9.285 1.460 9.790 1.800 ;
        RECT  7.955 3.345 8.415 3.625 ;
        RECT  8.185 1.255 8.415 3.625 ;
        RECT  7.950 3.395 8.290 3.680 ;
        RECT  9.930 0.910 10.310 1.250 ;
        RECT  9.780 2.620 10.310 2.960 ;
        RECT  10.025 0.910 10.310 2.960 ;
        RECT  9.555 2.675 9.840 3.870 ;
        RECT  9.550 3.510 9.840 3.870 ;
        RECT  4.890 3.105 6.90 3.135 ;
        RECT  4.890 3.105 6.30 3.335 ;
    END
END LSOGCPX0

MACRO LSOGCNX8
    CLASS CORE ;
    FOREIGN LSOGCNX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.380 1.105 18.720 3.740 ;
        RECT  17.765 2.250 18.720 2.590 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.590 3.470 11.300 3.850 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.795 2.250 16.515 2.650 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.869  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.060 2.660 3.400 4.180 ;
        RECT  3.060 1.015 3.400 1.355 ;
        RECT  3.060 1.015 3.310 4.180 ;
        RECT  1.615 2.005 3.310 2.350 ;
        RECT  1.615 1.030 1.960 4.180 ;
        RECT  1.385 1.640 1.960 2.295 ;
        RECT  0.180 1.955 1.960 2.295 ;
        RECT  0.180 1.045 0.520 4.215 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.631  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.430 2.040 9.325 2.630 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  17.660 2.820 18.000 5.280 ;
        RECT  16.175 2.885 16.515 5.280 ;
        RECT  13.755 3.515 14.095 5.280 ;
        RECT  12.335 3.530 12.675 5.280 ;
        RECT  9.575 2.750 9.915 5.280 ;
        RECT  7.135 2.560 7.480 5.280 ;
        RECT  4.780 2.560 5.120 5.280 ;
        RECT  3.780 2.660 4.120 5.280 ;
        RECT  2.340 2.660 2.680 5.280 ;
        RECT  0.900 2.645 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  17.660 -0.400 18.000 1.495 ;
        RECT  16.160 -0.400 16.500 1.250 ;
        RECT  13.780 -0.400 14.120 1.515 ;
        RECT  11.460 -0.400 11.800 1.580 ;
        RECT  10.060 -0.400 10.400 0.970 ;
        RECT  8.580 -0.400 8.925 1.340 ;
        RECT  7.140 -0.400 7.480 1.375 ;
        RECT  5.700 -0.400 6.040 1.375 ;
        RECT  3.780 -0.400 4.600 1.460 ;
        RECT  2.340 -0.400 2.680 1.385 ;
        RECT  0.900 -0.400 1.240 1.375 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  9.300 1.055 9.640 1.800 ;
        RECT  7.860 1.570 9.640 1.800 ;
        RECT  4.975 1.015 5.320 2.180 ;
        RECT  6.415 1.015 6.760 2.180 ;
        RECT  3.540 1.840 8.200 2.180 ;
        RECT  7.860 1.035 8.200 3.200 ;
        RECT  7.860 2.860 8.630 3.200 ;
        RECT  8.290 2.860 8.630 3.825 ;
        RECT  5.985 1.840 6.330 3.885 ;
        RECT  9.585 2.040 11.000 2.380 ;
        RECT  10.660 1.270 11.000 3.030 ;
        RECT  10.660 2.690 11.265 3.030 ;
        RECT  12.260 1.235 12.600 2.850 ;
        RECT  11.875 2.510 12.750 2.850 ;
        RECT  11.875 2.510 12.105 3.870 ;
        RECT  11.615 3.530 12.105 3.870 ;
        RECT  12.830 0.630 13.170 1.490 ;
        RECT  12.830 1.150 13.320 1.490 ;
        RECT  12.980 2.740 15.010 3.080 ;
        RECT  12.980 1.150 13.210 3.805 ;
        RECT  12.980 3.465 13.395 3.805 ;
        RECT  13.500 1.945 15.030 2.285 ;
        RECT  14.970 1.020 15.565 1.360 ;
        RECT  15.335 1.480 16.780 1.710 ;
        RECT  16.440 1.480 16.780 1.820 ;
        RECT  15.335 1.020 15.565 3.695 ;
        RECT  14.905 3.355 15.565 3.695 ;
        RECT  16.960 0.910 17.300 1.250 ;
        RECT  17.010 0.910 17.300 3.170 ;
        RECT  16.745 2.830 17.040 4.145 ;
        RECT  3.540 1.840 7.20 2.180 ;
        RECT  12.980 2.740 14.80 3.080 ;
    END
END LSOGCNX8

MACRO LSOGCNX6
    CLASS CORE ;
    FOREIGN LSOGCNX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.860 1.105 16.200 3.740 ;
        RECT  15.245 2.250 16.200 2.590 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.070 3.470 8.780 3.850 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.275 2.250 13.995 2.650 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.689  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.340 0.710 2.680 4.080 ;
        RECT  0.895 2.005 2.680 2.350 ;
        RECT  0.895 0.710 1.240 4.080 ;
        RECT  0.755 1.640 1.240 2.020 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.265  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.940 2.040 6.805 2.630 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.140 2.820 15.480 5.280 ;
        RECT  13.655 2.885 13.995 5.280 ;
        RECT  11.235 3.515 11.575 5.280 ;
        RECT  9.975 3.705 10.315 5.280 ;
        RECT  7.210 2.750 7.550 5.280 ;
        RECT  4.910 2.560 5.250 5.280 ;
        RECT  3.060 2.660 3.400 5.280 ;
        RECT  1.620 2.660 1.960 5.280 ;
        RECT  0.180 2.645 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.140 -0.400 15.480 1.495 ;
        RECT  13.640 -0.400 13.980 1.250 ;
        RECT  11.260 -0.400 11.600 1.515 ;
        RECT  8.940 -0.400 9.280 1.580 ;
        RECT  7.540 -0.400 7.880 0.970 ;
        RECT  6.060 -0.400 6.405 1.350 ;
        RECT  4.620 -0.400 4.960 1.495 ;
        RECT  3.100 -0.400 3.440 1.610 ;
        RECT  1.620 -0.400 1.960 1.620 ;
        RECT  0.180 -0.400 0.520 1.610 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  6.780 1.155 7.120 1.810 ;
        RECT  5.340 1.580 7.120 1.810 ;
        RECT  3.895 1.155 4.240 2.180 ;
        RECT  5.340 1.155 5.680 2.180 ;
        RECT  2.910 1.840 5.710 2.180 ;
        RECT  5.480 1.580 5.710 3.200 ;
        RECT  5.480 2.860 6.400 3.200 ;
        RECT  6.060 2.860 6.400 3.825 ;
        RECT  3.755 1.840 4.100 3.885 ;
        RECT  7.035 2.040 8.480 2.380 ;
        RECT  8.140 1.270 8.480 3.030 ;
        RECT  8.140 2.690 8.855 3.030 ;
        RECT  9.740 1.235 10.080 2.285 ;
        RECT  9.475 1.945 10.230 2.285 ;
        RECT  9.475 1.945 9.705 3.305 ;
        RECT  9.215 2.965 9.705 3.305 ;
        RECT  10.310 0.630 10.650 1.490 ;
        RECT  10.310 1.150 10.800 1.490 ;
        RECT  10.460 1.150 10.690 3.240 ;
        RECT  10.460 2.740 12.490 3.080 ;
        RECT  10.460 2.740 10.875 3.240 ;
        RECT  10.980 1.945 12.510 2.285 ;
        RECT  12.450 1.020 13.045 1.360 ;
        RECT  12.815 1.480 14.260 1.710 ;
        RECT  13.920 1.480 14.260 1.820 ;
        RECT  12.815 1.020 13.045 3.695 ;
        RECT  12.385 3.355 13.045 3.695 ;
        RECT  14.440 0.910 14.780 1.250 ;
        RECT  14.490 0.910 14.780 3.170 ;
        RECT  14.225 2.830 14.520 4.145 ;
        RECT  2.910 1.840 4.60 2.180 ;
        RECT  10.460 2.740 11.30 3.080 ;
    END
END LSOGCNX6

MACRO LSOGCNX4
    CLASS CORE ;
    FOREIGN LSOGCNX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 1.105 14.310 3.740 ;
        RECT  13.355 2.250 14.310 2.590 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.180 3.470 6.890 3.850 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.385 2.250 12.105 2.650 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 2.760 1.960 4.010 ;
        RECT  1.620 1.015 1.960 1.355 ;
        RECT  1.620 1.015 1.870 4.010 ;
        RECT  0.125 2.005 1.870 2.350 ;
        RECT  0.125 1.030 0.520 4.020 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.889  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.645 2.040 4.285 2.630 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.250 2.820 13.590 5.280 ;
        RECT  11.765 2.885 12.105 5.280 ;
        RECT  9.345 3.515 9.685 5.280 ;
        RECT  7.925 3.530 8.265 5.280 ;
        RECT  5.365 2.750 5.705 5.280 ;
        RECT  4.640 2.560 4.980 5.280 ;
        RECT  2.335 2.760 2.680 5.280 ;
        RECT  0.900 2.760 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.250 -0.400 13.590 1.495 ;
        RECT  11.750 -0.400 12.090 1.250 ;
        RECT  9.370 -0.400 9.710 1.515 ;
        RECT  6.820 -0.400 7.160 1.580 ;
        RECT  5.220 -0.400 5.560 1.395 ;
        RECT  3.780 -0.400 4.125 1.155 ;
        RECT  2.340 -0.400 2.680 1.340 ;
        RECT  0.900 -0.400 1.240 1.385 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  4.500 1.055 4.840 1.615 ;
        RECT  3.060 1.385 4.840 1.615 ;
        RECT  2.100 1.840 3.400 2.180 ;
        RECT  3.060 0.850 3.400 3.200 ;
        RECT  3.060 2.860 3.830 3.200 ;
        RECT  3.490 2.860 3.830 3.825 ;
        RECT  4.740 2.025 6.360 2.330 ;
        RECT  6.020 1.240 6.360 3.055 ;
        RECT  6.020 2.715 6.855 3.055 ;
        RECT  7.620 1.235 7.960 2.850 ;
        RECT  7.465 2.510 8.340 2.850 ;
        RECT  7.465 2.510 7.695 3.870 ;
        RECT  7.205 3.530 7.695 3.870 ;
        RECT  8.420 0.630 8.760 1.490 ;
        RECT  8.420 1.150 8.910 1.490 ;
        RECT  8.570 2.740 10.600 3.080 ;
        RECT  8.570 1.150 8.800 3.805 ;
        RECT  8.570 3.465 8.985 3.805 ;
        RECT  9.090 1.945 10.620 2.285 ;
        RECT  10.560 1.020 11.155 1.360 ;
        RECT  10.925 1.480 12.370 1.710 ;
        RECT  12.030 1.480 12.370 1.820 ;
        RECT  10.925 1.020 11.155 3.695 ;
        RECT  10.495 3.355 11.155 3.695 ;
        RECT  12.550 0.910 12.890 1.250 ;
        RECT  12.600 0.910 12.890 3.170 ;
        RECT  12.335 2.830 12.630 4.145 ;
        RECT  8.570 2.740 9.20 3.080 ;
    END
END LSOGCNX4

MACRO LSOGCNX3
    CLASS CORE ;
    FOREIGN LSOGCNX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.340 1.105 13.680 3.740 ;
        RECT  12.725 2.250 13.680 2.590 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.550 3.470 6.260 3.850 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.755 2.250 11.475 2.650 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.345  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 2.760 1.240 4.180 ;
        RECT  0.755 0.700 1.240 1.610 ;
        RECT  0.755 0.700 1.060 3.100 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.704  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.015 2.250 3.655 2.630 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.620 2.820 12.960 5.280 ;
        RECT  11.135 2.885 11.475 5.280 ;
        RECT  8.715 3.515 9.055 5.280 ;
        RECT  7.295 3.530 7.635 5.280 ;
        RECT  4.735 2.750 5.075 5.280 ;
        RECT  3.925 2.860 4.265 5.280 ;
        RECT  1.615 2.860 1.960 5.280 ;
        RECT  0.180 2.760 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.620 -0.400 12.960 1.495 ;
        RECT  11.120 -0.400 11.460 1.250 ;
        RECT  8.740 -0.400 9.080 1.515 ;
        RECT  6.140 -0.400 6.480 1.620 ;
        RECT  4.500 -0.400 4.840 1.395 ;
        RECT  3.060 -0.400 3.405 1.340 ;
        RECT  1.620 -0.400 1.960 1.340 ;
        RECT  0.180 -0.400 0.520 1.620 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.780 1.055 4.120 1.800 ;
        RECT  2.340 1.570 4.120 1.800 ;
        RECT  1.290 1.840 2.680 2.180 ;
        RECT  2.340 1.035 2.680 3.200 ;
        RECT  2.340 2.860 3.115 3.200 ;
        RECT  2.775 2.860 3.115 3.825 ;
        RECT  3.955 2.030 5.680 2.365 ;
        RECT  5.305 1.280 5.680 3.055 ;
        RECT  5.305 2.715 6.225 3.055 ;
        RECT  6.940 1.275 7.280 2.850 ;
        RECT  6.835 2.510 7.710 2.850 ;
        RECT  6.835 2.510 7.065 3.870 ;
        RECT  6.575 3.530 7.065 3.870 ;
        RECT  7.790 0.630 8.130 1.490 ;
        RECT  7.790 1.150 8.280 1.490 ;
        RECT  7.940 2.740 9.970 3.080 ;
        RECT  7.940 1.150 8.170 3.805 ;
        RECT  7.940 3.465 8.355 3.805 ;
        RECT  8.460 1.945 9.990 2.285 ;
        RECT  9.930 1.020 10.525 1.360 ;
        RECT  10.295 1.480 11.740 1.710 ;
        RECT  11.400 1.480 11.740 1.820 ;
        RECT  10.295 1.020 10.525 3.695 ;
        RECT  9.865 3.355 10.525 3.695 ;
        RECT  11.920 0.910 12.260 1.250 ;
        RECT  11.970 0.910 12.260 3.170 ;
        RECT  11.705 2.830 12.000 4.145 ;
        RECT  7.940 2.740 8.50 3.080 ;
    END
END LSOGCNX3

MACRO LSOGCNX2
    CLASS CORE ;
    FOREIGN LSOGCNX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 1.105 12.420 3.740 ;
        RECT  11.465 2.250 12.420 2.590 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.290 3.470 5.000 3.850 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.495 2.250 10.215 2.650 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.901  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.160 1.245 3.500 ;
        RECT  0.755 1.015 1.240 1.355 ;
        RECT  0.755 2.250 1.135 3.500 ;
        RECT  0.755 1.015 0.985 3.500 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.518  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.655 2.395 3.025 3.240 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.360 2.820 11.700 5.280 ;
        RECT  9.875 2.885 10.215 5.280 ;
        RECT  7.455 3.515 7.795 5.280 ;
        RECT  6.035 3.530 6.375 5.280 ;
        RECT  3.475 2.750 3.815 5.280 ;
        RECT  1.625 3.150 1.965 5.280 ;
        RECT  0.180 2.790 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.360 -0.400 11.700 1.495 ;
        RECT  9.860 -0.400 10.200 1.250 ;
        RECT  7.480 -0.400 7.820 1.515 ;
        RECT  4.880 -0.400 5.220 1.620 ;
        RECT  3.130 -0.400 3.470 1.395 ;
        RECT  1.620 -0.400 1.960 1.235 ;
        RECT  0.180 -0.400 0.520 1.365 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.450 1.465 2.680 1.695 ;
        RECT  2.340 1.135 2.680 1.695 ;
        RECT  1.290 1.695 1.680 2.035 ;
        RECT  1.450 1.465 1.680 2.835 ;
        RECT  1.450 2.605 2.425 2.835 ;
        RECT  2.195 2.605 2.425 3.760 ;
        RECT  2.195 3.470 3.115 3.760 ;
        RECT  4.045 1.280 4.420 1.620 ;
        RECT  2.010 1.925 4.275 2.165 ;
        RECT  2.010 1.925 2.350 2.220 ;
        RECT  4.045 1.280 4.275 2.925 ;
        RECT  4.045 2.585 4.965 2.925 ;
        RECT  5.680 1.275 6.020 2.850 ;
        RECT  5.575 2.510 6.450 2.850 ;
        RECT  5.575 2.510 5.805 3.870 ;
        RECT  5.315 3.530 5.805 3.870 ;
        RECT  6.530 0.630 6.870 1.490 ;
        RECT  6.530 1.150 7.020 1.490 ;
        RECT  6.680 2.740 8.710 3.080 ;
        RECT  6.680 1.150 6.910 3.805 ;
        RECT  6.680 3.465 7.095 3.805 ;
        RECT  7.200 1.945 8.730 2.285 ;
        RECT  8.670 1.020 9.265 1.360 ;
        RECT  9.035 1.480 10.480 1.710 ;
        RECT  10.140 1.480 10.480 1.820 ;
        RECT  9.035 1.020 9.265 3.695 ;
        RECT  8.605 3.355 9.265 3.695 ;
        RECT  10.660 0.910 11.000 1.250 ;
        RECT  10.710 0.910 11.000 3.170 ;
        RECT  10.445 2.830 10.740 4.145 ;
        RECT  2.010 1.925 3.00 2.165 ;
        RECT  6.680 2.740 7.40 3.080 ;
    END
END LSOGCNX2

MACRO LSOGCNX1
    CLASS CORE ;
    FOREIGN LSOGCNX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 0.820 10.585 4.180 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.110 3.460 3.720 3.860 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 2.250 8.280 2.655 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.640 0.520 3.560 ;
        RECT  0.125 1.185 0.520 1.525 ;
        RECT  0.125 1.185 0.355 3.560 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.333  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.840 2.250 2.405 2.685 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 3.610 9.810 5.280 ;
        RECT  8.015 3.850 8.355 5.280 ;
        RECT  5.995 3.400 6.335 5.280 ;
        RECT  4.735 3.530 5.075 5.280 ;
        RECT  2.470 2.920 2.810 5.280 ;
        RECT  0.740 3.960 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.430 -0.400 9.770 0.915 ;
        RECT  8.130 -0.400 8.470 0.905 ;
        RECT  5.700 -0.400 6.040 0.970 ;
        RECT  3.540 -0.400 3.880 0.995 ;
        RECT  2.340 -0.400 2.680 0.995 ;
        RECT  0.940 -0.400 1.280 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.800 1.275 1.880 1.560 ;
        RECT  0.590 1.825 1.030 2.165 ;
        RECT  0.800 1.275 1.030 3.155 ;
        RECT  0.800 2.925 1.700 3.155 ;
        RECT  1.470 2.925 1.700 4.215 ;
        RECT  1.470 3.875 2.110 4.215 ;
        RECT  2.940 1.305 3.280 2.020 ;
        RECT  1.260 1.790 3.850 2.020 ;
        RECT  1.260 1.790 1.600 2.215 ;
        RECT  3.620 1.790 3.850 2.980 ;
        RECT  3.620 2.640 3.960 2.980 ;
        RECT  4.400 1.300 4.740 2.165 ;
        RECT  4.190 1.825 4.860 2.165 ;
        RECT  4.190 1.825 4.420 3.955 ;
        RECT  3.950 3.615 4.420 3.955 ;
        RECT  6.650 0.785 6.980 1.115 ;
        RECT  6.650 0.785 6.970 1.125 ;
        RECT  6.650 0.785 6.880 2.035 ;
        RECT  5.550 1.805 6.880 2.035 ;
        RECT  5.550 1.805 5.890 2.145 ;
        RECT  4.965 0.630 5.440 0.970 ;
        RECT  5.090 0.630 5.440 1.600 ;
        RECT  5.090 0.630 5.425 1.610 ;
        RECT  5.090 0.630 5.320 2.680 ;
        RECT  6.650 2.310 6.990 2.680 ;
        RECT  5.090 2.450 6.990 2.680 ;
        RECT  5.295 2.450 5.635 3.065 ;
        RECT  7.140 1.285 7.480 1.625 ;
        RECT  7.220 1.285 7.480 2.020 ;
        RECT  7.220 1.790 8.990 2.020 ;
        RECT  8.650 1.790 8.990 2.145 ;
        RECT  7.220 1.285 7.450 4.250 ;
        RECT  7.185 3.910 7.525 4.250 ;
        RECT  8.930 1.275 9.535 1.560 ;
        RECT  9.305 1.275 9.535 3.220 ;
        RECT  8.585 2.880 9.535 3.220 ;
        RECT  8.585 2.880 8.925 4.140 ;
        RECT  1.260 1.790 2.60 2.020 ;
    END
END LSOGCNX1

MACRO LSOGCNX0
    CLASS CORE ;
    FOREIGN LSOGCNX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CGOBS
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.569  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.500 2.250 9.955 2.980 ;
        RECT  9.500 1.170 9.890 1.510 ;
        RECT  9.500 1.170 9.730 2.980 ;
        END
    END CGOBS
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.610 1.640 4.285 2.020 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.315 2.175 8.695 2.600 ;
        RECT  7.800 2.175 8.695 2.405 ;
        RECT  7.800 1.570 8.030 2.405 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.640 0.520 3.240 ;
        RECT  0.125 1.150 0.520 1.490 ;
        RECT  0.125 1.150 0.355 3.240 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.540 2.405 2.165 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.445 3.590 9.785 5.280 ;
        RECT  7.770 3.555 8.130 5.280 ;
        RECT  4.775 3.510 5.715 5.280 ;
        RECT  5.375 3.340 5.715 5.280 ;
        RECT  2.210 3.405 2.550 5.280 ;
        RECT  0.980 2.450 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  9.550 -0.400 9.890 0.710 ;
        RECT  8.150 -0.400 8.490 0.710 ;
        RECT  6.700 -0.400 6.930 1.210 ;
        RECT  5.875 1.340 6.895 1.630 ;
        RECT  6.655 1.065 6.895 1.630 ;
        RECT  3.980 -0.400 5.085 0.870 ;
        RECT  3.980 -0.400 4.320 1.365 ;
        RECT  2.380 -0.400 2.720 1.310 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.555 1.025 1.920 1.310 ;
        RECT  1.555 1.025 1.900 1.340 ;
        RECT  0.630 1.815 0.970 2.155 ;
        RECT  0.630 1.925 1.785 2.155 ;
        RECT  1.555 1.025 1.785 2.715 ;
        RECT  1.555 2.430 2.550 2.715 ;
        RECT  3.150 1.025 3.520 1.365 ;
        RECT  3.150 2.530 3.780 2.870 ;
        RECT  3.150 1.025 3.380 3.175 ;
        RECT  1.550 2.945 3.380 3.175 ;
        RECT  1.550 2.945 1.840 3.660 ;
        RECT  4.800 1.245 5.085 3.270 ;
        RECT  3.975 3.040 5.085 3.270 ;
        RECT  3.975 3.040 4.315 3.570 ;
        RECT  5.315 0.630 6.470 0.915 ;
        RECT  5.315 0.630 5.545 2.965 ;
        RECT  5.315 2.625 6.835 2.965 ;
        RECT  6.495 2.625 6.835 3.155 ;
        RECT  6.495 2.625 6.780 3.160 ;
        RECT  5.775 1.860 6.060 2.200 ;
        RECT  5.775 1.970 7.110 2.200 ;
        RECT  6.825 1.970 7.110 2.310 ;
        RECT  7.310 1.110 8.490 1.340 ;
        RECT  8.260 1.110 8.490 1.870 ;
        RECT  7.125 1.340 7.570 1.680 ;
        RECT  8.260 1.580 8.810 1.870 ;
        RECT  7.340 1.110 7.570 3.060 ;
        RECT  7.310 2.830 7.540 3.640 ;
        RECT  6.830 3.385 7.540 3.640 ;
        RECT  6.815 3.410 7.155 3.695 ;
        RECT  8.750 1.060 9.270 1.350 ;
        RECT  9.040 1.060 9.270 3.115 ;
        RECT  8.365 2.830 9.270 3.115 ;
        RECT  8.365 2.830 8.985 3.170 ;
        RECT  8.365 2.830 8.705 4.130 ;
    END
END LSOGCNX0

MACRO LSGCPX8
    CLASS CORE ;
    FOREIGN LSGCPX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.470 3.660 3.985 ;
        RECT  3.260 3.325 3.535 3.985 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.147  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.595 0.720 14.995 4.180 ;
        RECT  11.755 1.965 14.995 2.305 ;
        RECT  13.155 0.720 13.495 4.180 ;
        RECT  11.715 2.705 12.105 4.195 ;
        RECT  11.755 0.725 12.105 4.195 ;
        RECT  11.715 0.725 12.105 1.700 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.205 1.640 6.805 2.240 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.445 4.915 2.020 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.875 -0.400 14.215 1.700 ;
        RECT  12.435 -0.400 12.775 1.710 ;
        RECT  10.995 -0.400 11.340 1.555 ;
        RECT  8.695 -0.400 9.035 1.515 ;
        RECT  6.395 -0.400 6.735 1.410 ;
        RECT  4.750 -0.400 5.090 0.920 ;
        RECT  3.140 -0.400 3.490 1.320 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  13.875 2.705 14.215 5.280 ;
        RECT  12.430 2.705 12.775 5.280 ;
        RECT  10.995 2.660 11.345 5.280 ;
        RECT  9.555 2.770 9.895 5.280 ;
        RECT  8.115 2.770 8.455 5.280 ;
        RECT  6.675 2.915 7.015 5.280 ;
        RECT  4.785 3.910 5.125 5.280 ;
        RECT  2.730 2.615 3.380 2.955 ;
        RECT  2.730 2.615 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.320 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  0.240 0.830 0.580 1.170 ;
        RECT  0.240 0.940 2.320 1.170 ;
        RECT  1.715 0.940 2.320 1.320 ;
        RECT  1.715 0.940 1.945 3.085 ;
        RECT  1.715 2.725 2.230 3.085 ;
        RECT  1.255 2.855 2.230 3.085 ;
        RECT  1.255 2.855 1.540 4.210 ;
        RECT  3.950 1.090 4.305 1.880 ;
        RECT  2.965 1.565 4.305 1.880 ;
        RECT  4.075 1.090 4.305 2.480 ;
        RECT  4.210 2.250 4.550 2.815 ;
        RECT  5.320 0.630 5.890 0.970 ;
        RECT  5.320 0.630 5.550 1.370 ;
        RECT  2.175 2.000 2.470 2.340 ;
        RECT  5.145 1.145 5.375 2.480 ;
        RECT  2.175 2.110 3.840 2.340 ;
        RECT  3.610 2.110 3.840 2.940 ;
        RECT  3.750 2.710 3.980 3.210 ;
        RECT  4.835 2.250 5.165 3.525 ;
        RECT  3.785 3.045 5.165 3.275 ;
        RECT  4.825 3.045 5.165 3.525 ;
        RECT  5.645 1.580 5.935 3.245 ;
        RECT  5.395 2.905 5.935 3.245 ;
        RECT  5.395 2.910 6.255 3.245 ;
        RECT  7.545 1.175 7.890 2.405 ;
        RECT  9.845 1.175 10.185 2.405 ;
        RECT  7.395 2.065 11.525 2.405 ;
        RECT  8.830 2.065 9.175 3.870 ;
        RECT  7.395 2.065 7.735 3.880 ;
        RECT  10.275 2.065 10.615 3.880 ;
        RECT  0.240 0.940 1.50 1.170 ;
        RECT  7.395 2.065 10.10 2.405 ;
    END
END LSGCPX8

MACRO LSGCPX6
    CLASS CORE ;
    FOREIGN LSGCPX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.415 3.660 3.985 ;
        RECT  3.275 3.325 3.615 3.985 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.689  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.250 0.790 13.590 4.080 ;
        RECT  11.850 2.250 13.590 2.630 ;
        RECT  11.810 2.660 12.150 4.080 ;
        RECT  11.850 0.790 12.150 4.080 ;
        RECT  11.810 0.790 12.150 1.700 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.365 2.150 6.870 2.650 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.610 5.035 2.020 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.970 -0.400 14.310 1.700 ;
        RECT  12.530 -0.400 12.870 1.700 ;
        RECT  11.090 -0.400 11.430 1.435 ;
        RECT  8.785 -0.400 9.130 1.495 ;
        RECT  6.340 -0.400 6.680 0.950 ;
        RECT  4.840 -0.400 5.180 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.970 2.660 14.310 5.280 ;
        RECT  12.530 2.860 12.870 5.280 ;
        RECT  11.090 2.960 11.430 5.280 ;
        RECT  9.650 2.960 9.995 5.280 ;
        RECT  8.210 2.960 8.550 5.280 ;
        RECT  6.765 2.960 7.110 5.280 ;
        RECT  5.335 3.440 5.675 5.280 ;
        RECT  2.745 2.615 3.380 2.955 ;
        RECT  2.745 2.615 3.045 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.320 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  0.240 0.830 0.580 1.170 ;
        RECT  0.240 0.940 2.350 1.170 ;
        RECT  1.715 0.940 2.350 1.320 ;
        RECT  1.715 0.940 1.945 3.085 ;
        RECT  1.715 2.725 2.230 3.085 ;
        RECT  1.255 2.855 2.230 3.085 ;
        RECT  1.255 2.855 1.540 4.210 ;
        RECT  4.040 1.090 4.380 1.440 ;
        RECT  4.040 1.090 4.305 1.880 ;
        RECT  2.965 1.565 4.305 1.880 ;
        RECT  4.075 1.090 4.305 2.480 ;
        RECT  4.305 2.250 4.645 2.815 ;
        RECT  5.410 0.630 5.980 0.970 ;
        RECT  5.410 0.630 5.640 1.430 ;
        RECT  2.175 2.000 2.470 2.340 ;
        RECT  2.175 2.110 3.840 2.340 ;
        RECT  3.610 2.110 3.840 2.940 ;
        RECT  3.610 2.710 4.075 2.940 ;
        RECT  3.845 2.710 4.075 3.275 ;
        RECT  5.265 1.200 5.495 3.210 ;
        RECT  4.875 2.980 5.495 3.210 ;
        RECT  3.845 3.045 5.105 3.275 ;
        RECT  4.605 3.045 5.105 3.820 ;
        RECT  5.895 1.410 6.685 1.750 ;
        RECT  5.895 1.410 6.125 2.110 ;
        RECT  5.755 1.880 6.095 3.175 ;
        RECT  6.055 2.945 6.395 3.780 ;
        RECT  7.640 1.185 7.980 2.250 ;
        RECT  9.940 1.190 10.280 2.250 ;
        RECT  7.490 1.910 11.620 2.250 ;
        RECT  7.490 1.910 7.830 3.880 ;
        RECT  8.930 1.910 9.270 3.880 ;
        RECT  10.370 1.910 10.710 3.880 ;
        RECT  0.240 0.940 1.40 1.170 ;
        RECT  7.490 1.910 10.60 2.250 ;
    END
END LSGCPX6

MACRO LSGCPX4
    CLASS CORE ;
    FOREIGN LSGCPX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.480 3.660 3.985 ;
        RECT  3.260 3.325 3.535 3.985 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.373  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.915 1.115 12.255 4.180 ;
        RECT  10.515 2.250 12.255 2.630 ;
        RECT  10.450 2.770 10.855 4.180 ;
        RECT  10.515 2.250 10.855 4.180 ;
        RECT  10.515 1.115 10.815 4.180 ;
        RECT  10.475 1.115 10.815 1.455 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.360 2.070 6.805 2.650 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.610 5.035 2.020 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.195 -0.400 11.535 1.455 ;
        RECT  9.755 -0.400 10.095 1.435 ;
        RECT  7.450 -0.400 7.795 1.420 ;
        RECT  4.840 -0.400 5.180 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.195 2.930 11.535 5.280 ;
        RECT  9.755 2.960 10.095 5.280 ;
        RECT  8.195 3.220 8.540 5.280 ;
        RECT  6.755 3.245 7.095 5.280 ;
        RECT  5.335 3.415 5.675 5.280 ;
        RECT  2.730 2.615 3.380 2.955 ;
        RECT  2.730 2.615 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.320 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  0.240 0.830 0.580 1.170 ;
        RECT  0.240 0.940 2.350 1.170 ;
        RECT  1.715 0.940 2.350 1.320 ;
        RECT  1.715 0.940 1.945 3.085 ;
        RECT  1.715 2.725 2.230 3.085 ;
        RECT  1.255 2.855 2.230 3.085 ;
        RECT  1.255 2.855 1.540 4.210 ;
        RECT  4.040 1.090 4.380 1.440 ;
        RECT  4.040 1.090 4.305 1.880 ;
        RECT  2.965 1.565 4.305 1.880 ;
        RECT  4.075 1.090 4.305 2.480 ;
        RECT  4.210 2.250 4.550 2.815 ;
        RECT  5.410 0.630 5.980 0.970 ;
        RECT  5.410 0.630 5.640 1.430 ;
        RECT  2.175 2.000 2.470 2.340 ;
        RECT  2.175 2.110 3.840 2.340 ;
        RECT  3.610 2.110 3.840 2.940 ;
        RECT  3.750 2.710 3.980 3.210 ;
        RECT  5.265 1.200 5.495 3.135 ;
        RECT  4.780 2.905 5.495 3.135 ;
        RECT  3.775 3.045 5.010 3.275 ;
        RECT  4.605 3.045 5.010 3.820 ;
        RECT  6.655 1.180 6.995 1.520 ;
        RECT  5.895 1.200 6.995 1.520 ;
        RECT  5.725 1.880 6.125 2.220 ;
        RECT  5.890 1.880 6.125 3.175 ;
        RECT  5.895 1.200 6.125 3.175 ;
        RECT  6.055 2.945 6.395 3.740 ;
        RECT  8.605 1.140 8.945 2.250 ;
        RECT  7.475 1.910 10.285 2.250 ;
        RECT  7.475 1.910 7.815 3.530 ;
        RECT  8.915 1.910 9.255 3.530 ;
        RECT  0.240 0.940 1.40 1.170 ;
        RECT  7.475 1.910 9.80 2.250 ;
    END
END LSGCPX4

MACRO LSGCPX3
    CLASS CORE ;
    FOREIGN LSGCPX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.480 3.660 3.985 ;
        RECT  3.260 3.325 3.535 3.985 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.345  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.515 2.250 11.215 2.630 ;
        RECT  10.450 2.760 10.855 4.180 ;
        RECT  10.515 2.250 10.855 4.180 ;
        RECT  10.515 0.790 10.815 4.180 ;
        RECT  10.475 0.790 10.815 1.695 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.635  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.360 2.070 6.805 2.650 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.610 5.035 2.020 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  11.195 -0.400 11.535 1.700 ;
        RECT  9.755 -0.400 10.095 1.435 ;
        RECT  7.450 -0.400 7.795 1.385 ;
        RECT  4.840 -0.400 5.180 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.195 2.860 11.535 5.280 ;
        RECT  9.755 3.130 10.095 5.280 ;
        RECT  8.195 3.130 8.540 5.280 ;
        RECT  6.755 3.135 7.095 5.280 ;
        RECT  5.335 3.415 5.675 5.280 ;
        RECT  2.730 2.615 3.380 2.955 ;
        RECT  2.730 2.615 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.320 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  0.240 0.830 0.580 1.170 ;
        RECT  0.240 0.940 2.350 1.170 ;
        RECT  1.715 0.940 2.350 1.320 ;
        RECT  1.715 0.940 1.945 3.085 ;
        RECT  1.715 2.725 2.230 3.085 ;
        RECT  1.255 2.855 2.230 3.085 ;
        RECT  1.255 2.855 1.540 4.210 ;
        RECT  4.040 1.090 4.380 1.440 ;
        RECT  4.040 1.090 4.305 1.880 ;
        RECT  2.965 1.565 4.305 1.880 ;
        RECT  4.075 1.090 4.305 2.480 ;
        RECT  4.210 2.250 4.550 2.815 ;
        RECT  5.410 0.630 5.980 0.970 ;
        RECT  5.410 0.630 5.640 1.430 ;
        RECT  2.175 2.000 2.470 2.340 ;
        RECT  2.175 2.110 3.840 2.340 ;
        RECT  3.610 2.110 3.840 2.940 ;
        RECT  3.750 2.710 3.980 3.220 ;
        RECT  5.265 1.200 5.495 3.135 ;
        RECT  4.780 2.905 5.495 3.135 ;
        RECT  3.770 3.045 5.010 3.275 ;
        RECT  4.605 3.045 5.010 3.820 ;
        RECT  6.655 1.180 6.995 1.520 ;
        RECT  5.895 1.200 6.995 1.520 ;
        RECT  5.725 1.880 6.125 3.175 ;
        RECT  5.895 1.200 6.125 3.175 ;
        RECT  6.055 2.945 6.395 3.740 ;
        RECT  8.605 1.080 8.945 2.220 ;
        RECT  7.475 1.880 10.285 2.220 ;
        RECT  8.915 1.880 9.255 3.435 ;
        RECT  7.475 1.880 7.815 3.450 ;
        RECT  0.240 0.940 1.40 1.170 ;
        RECT  7.475 1.880 9.40 2.220 ;
    END
END LSGCPX3

MACRO LSGCPX2
    CLASS CORE ;
    FOREIGN LSGCPX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.230 3.480 3.655 3.985 ;
        RECT  3.230 3.330 3.535 3.985 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 2.850 9.335 3.770 ;
        RECT  9.090 1.240 9.335 3.770 ;
        RECT  8.930 1.240 9.335 1.580 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.360 2.070 6.805 2.630 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.610 5.035 2.020 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  9.490 -0.400 9.830 0.710 ;
        RECT  8.360 -0.400 8.710 0.720 ;
        RECT  6.565 1.330 6.980 1.670 ;
        RECT  6.565 -0.400 6.910 1.670 ;
        RECT  4.840 -0.400 5.180 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.490 4.170 9.830 5.280 ;
        RECT  8.210 3.130 8.550 5.280 ;
        RECT  6.770 3.535 7.115 5.280 ;
        RECT  5.670 3.650 6.010 5.280 ;
        RECT  2.700 2.615 3.380 2.955 ;
        RECT  2.700 2.615 3.000 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.320 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  0.240 0.830 0.580 1.170 ;
        RECT  0.240 0.940 2.350 1.170 ;
        RECT  1.715 0.940 2.350 1.320 ;
        RECT  1.715 0.940 1.945 3.085 ;
        RECT  1.715 2.725 2.230 3.085 ;
        RECT  1.255 2.855 2.230 3.085 ;
        RECT  1.255 2.855 1.540 4.210 ;
        RECT  4.040 1.090 4.380 1.440 ;
        RECT  4.040 1.090 4.305 1.880 ;
        RECT  2.965 1.565 4.305 1.880 ;
        RECT  4.075 1.090 4.305 2.480 ;
        RECT  4.210 2.250 4.550 2.815 ;
        RECT  5.410 0.630 5.980 0.970 ;
        RECT  5.410 0.630 5.640 1.430 ;
        RECT  2.175 2.000 2.470 2.340 ;
        RECT  2.175 2.110 3.840 2.340 ;
        RECT  3.610 2.110 3.840 2.940 ;
        RECT  3.750 2.710 3.980 3.245 ;
        RECT  5.265 1.200 5.495 3.275 ;
        RECT  4.910 2.905 5.495 3.275 ;
        RECT  3.765 3.045 5.495 3.275 ;
        RECT  5.870 1.315 6.180 1.670 ;
        RECT  5.870 1.315 6.125 3.175 ;
        RECT  5.725 1.880 6.125 3.175 ;
        RECT  5.725 2.860 6.585 3.175 ;
        RECT  7.140 0.640 7.830 0.980 ;
        RECT  7.490 1.880 8.860 2.220 ;
        RECT  7.490 0.640 7.830 3.800 ;
        RECT  0.240 0.940 1.30 1.170 ;
    END
END LSGCPX2

MACRO LSGCPX1
    CLASS CORE ;
    FOREIGN LSGCPX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.505 3.660 3.985 ;
        RECT  3.260 3.480 3.645 3.985 ;
        RECT  3.260 3.360 3.535 3.985 ;
        RECT  3.260 3.325 3.520 3.985 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 2.860 9.335 4.180 ;
        RECT  9.090 1.240 9.335 4.180 ;
        RECT  8.930 1.240 9.335 1.580 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.311  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.360 2.070 6.805 2.630 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.610 5.035 2.020 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.360 -0.400 8.710 0.720 ;
        RECT  6.635 -0.400 6.980 1.670 ;
        RECT  4.840 -0.400 5.180 0.970 ;
        RECT  3.240 -0.400 3.580 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.210 3.540 8.550 5.280 ;
        RECT  6.770 3.535 7.115 5.280 ;
        RECT  5.670 3.650 6.010 5.280 ;
        RECT  2.730 2.615 3.380 2.955 ;
        RECT  2.730 2.615 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.320 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  0.240 0.830 0.580 1.170 ;
        RECT  0.240 0.940 2.350 1.170 ;
        RECT  1.715 0.940 2.350 1.320 ;
        RECT  1.715 0.940 1.945 3.085 ;
        RECT  1.715 2.725 2.230 3.085 ;
        RECT  1.255 2.855 2.230 3.085 ;
        RECT  1.255 2.855 1.540 4.210 ;
        RECT  4.040 1.090 4.380 1.440 ;
        RECT  4.040 1.090 4.305 1.880 ;
        RECT  2.965 1.565 4.305 1.880 ;
        RECT  4.075 1.090 4.305 2.480 ;
        RECT  4.210 2.250 4.550 2.815 ;
        RECT  5.410 0.630 5.980 0.970 ;
        RECT  5.410 0.630 5.640 1.430 ;
        RECT  2.175 2.000 2.470 2.340 ;
        RECT  2.175 2.110 3.840 2.340 ;
        RECT  3.610 2.110 3.840 2.940 ;
        RECT  3.750 2.710 3.980 3.275 ;
        RECT  5.265 1.200 5.495 3.275 ;
        RECT  4.910 2.905 5.495 3.275 ;
        RECT  3.750 3.045 5.495 3.275 ;
        RECT  5.870 1.315 6.180 1.670 ;
        RECT  5.870 1.315 6.125 2.110 ;
        RECT  5.725 1.880 6.010 3.175 ;
        RECT  5.725 2.860 6.585 3.175 ;
        RECT  7.340 0.640 7.900 0.980 ;
        RECT  7.670 1.880 8.860 2.220 ;
        RECT  7.670 0.640 7.900 3.800 ;
        RECT  7.490 3.460 7.900 3.800 ;
        RECT  0.240 0.940 1.20 1.170 ;
    END
END LSGCPX1

MACRO LSGCPX0
    CLASS CORE ;
    FOREIGN LSGCPX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.105 6.995 2.630 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.640 8.065 2.385 ;
        END
    END SE
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.640 0.520 3.240 ;
        RECT  0.125 1.150 0.520 1.490 ;
        RECT  0.125 1.150 0.355 3.240 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.535 2.405 2.160 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.500 -0.400 7.840 0.655 ;
        RECT  6.300 -0.400 6.640 0.655 ;
        RECT  4.095 1.340 4.705 1.680 ;
        RECT  4.475 -0.400 4.705 1.680 ;
        RECT  2.610 -0.400 3.405 0.715 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.300 4.015 8.640 5.280 ;
        RECT  6.635 3.700 6.975 5.280 ;
        RECT  3.925 3.100 4.265 5.280 ;
        RECT  2.620 3.750 2.960 5.280 ;
        RECT  0.980 2.640 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.555 0.630 2.150 0.945 ;
        RECT  0.630 1.815 0.970 2.155 ;
        RECT  0.630 1.925 1.785 2.155 ;
        RECT  1.555 0.630 1.785 2.985 ;
        RECT  1.555 2.645 2.120 2.985 ;
        RECT  2.765 1.275 3.405 1.615 ;
        RECT  2.765 1.275 3.090 2.250 ;
        RECT  2.765 1.275 3.050 3.520 ;
        RECT  1.780 3.290 3.050 3.520 ;
        RECT  1.780 3.290 2.120 3.685 ;
        RECT  3.635 0.640 4.245 0.980 ;
        RECT  3.635 0.640 3.865 2.855 ;
        RECT  4.875 2.385 5.215 2.855 ;
        RECT  3.280 2.570 5.215 2.855 ;
        RECT  3.280 2.570 3.565 3.155 ;
        RECT  5.395 1.345 5.735 1.680 ;
        RECT  5.505 1.345 5.735 4.095 ;
        RECT  5.325 3.545 5.735 4.095 ;
        RECT  5.325 3.755 6.185 4.095 ;
        RECT  5.965 1.345 7.455 1.635 ;
        RECT  5.965 1.345 6.255 1.910 ;
        RECT  7.225 1.345 7.455 3.200 ;
        RECT  7.225 2.860 8.010 3.200 ;
        RECT  4.935 0.885 8.705 1.115 ;
        RECT  8.300 0.885 8.705 1.390 ;
        RECT  4.935 0.885 5.165 2.145 ;
        RECT  4.205 1.910 5.165 2.145 ;
        RECT  4.205 1.910 4.545 2.150 ;
        RECT  8.475 0.885 8.705 3.785 ;
        RECT  7.500 3.555 8.705 3.785 ;
        RECT  7.500 3.555 7.840 3.970 ;
        RECT  4.935 0.885 7.80 1.115 ;
    END
END LSGCPX0

MACRO LSGCNX8
    CLASS CORE ;
    FOREIGN LSGCNX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.295 3.665 3.895 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 3.310 4.330 3.880 ;
        END
    END SE
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.633  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.525 1.800 7.285 2.140 ;
        RECT  6.425 2.225 6.805 2.630 ;
        RECT  6.525 1.800 6.805 2.630 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.857  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.715 2.035 14.995 2.335 ;
        RECT  14.595 0.700 14.995 2.335 ;
        RECT  13.875 2.035 14.215 3.770 ;
        RECT  13.155 0.700 13.495 2.335 ;
        RECT  12.555 2.035 12.895 3.770 ;
        RECT  11.235 2.745 12.055 3.085 ;
        RECT  11.715 1.130 12.055 3.085 ;
        RECT  11.235 2.745 11.575 3.770 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.875 -0.400 14.215 1.700 ;
        RECT  12.435 -0.400 12.775 1.805 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  9.675 -0.400 10.015 1.295 ;
        RECT  8.235 -0.400 8.575 1.390 ;
        RECT  6.795 -0.400 7.135 1.390 ;
        RECT  5.090 -0.400 5.320 0.970 ;
        RECT  3.195 -0.400 3.480 1.320 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.595 2.735 14.935 5.280 ;
        RECT  13.315 4.170 13.655 5.280 ;
        RECT  11.995 4.170 12.335 5.280 ;
        RECT  10.675 4.170 11.015 5.280 ;
        RECT  8.335 2.840 8.675 5.280 ;
        RECT  5.395 3.570 6.205 5.280 ;
        RECT  2.730 2.670 3.380 3.010 ;
        RECT  2.730 2.670 3.030 5.280 ;
        RECT  0.740 2.720 1.045 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.505 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  1.275 2.120 1.505 4.210 ;
        RECT  1.275 3.870 2.040 4.210 ;
        RECT  0.180 0.830 0.520 1.170 ;
        RECT  0.180 0.940 2.345 1.170 ;
        RECT  1.735 0.940 2.345 1.280 ;
        RECT  1.735 0.940 1.965 3.065 ;
        RECT  1.735 2.725 2.230 3.065 ;
        RECT  4.170 1.090 4.400 2.350 ;
        RECT  2.870 2.010 4.550 2.350 ;
        RECT  4.210 2.010 4.550 3.010 ;
        RECT  3.710 0.630 4.860 0.860 ;
        RECT  5.550 0.630 6.185 0.950 ;
        RECT  4.630 0.630 4.860 1.430 ;
        RECT  5.550 0.630 5.780 1.430 ;
        RECT  4.630 1.200 5.780 1.430 ;
        RECT  3.710 0.630 3.940 1.780 ;
        RECT  2.195 1.550 3.940 1.780 ;
        RECT  2.195 1.510 2.535 1.850 ;
        RECT  4.780 1.200 5.010 3.780 ;
        RECT  4.635 3.440 5.010 3.780 ;
        RECT  6.010 1.310 6.295 1.960 ;
        RECT  5.240 1.660 6.295 1.960 ;
        RECT  5.240 1.660 5.605 2.970 ;
        RECT  8.955 0.955 9.295 2.610 ;
        RECT  10.395 0.955 10.735 2.490 ;
        RECT  7.515 1.050 7.855 2.610 ;
        RECT  7.515 2.270 11.335 2.490 ;
        RECT  8.955 2.150 11.335 2.490 ;
        RECT  7.185 2.370 9.825 2.610 ;
        RECT  7.185 2.370 7.525 3.880 ;
        RECT  9.485 2.150 9.825 3.880 ;
        RECT  0.180 0.940 1.80 1.170 ;
        RECT  7.515 2.270 10.80 2.490 ;
        RECT  8.955 2.150 10.30 2.490 ;
        RECT  7.185 2.370 8.70 2.610 ;
    END
END LSGCNX8

MACRO LSGCNX6
    CLASS CORE ;
    FOREIGN LSGCNX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.295 3.665 3.895 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 3.310 4.330 3.880 ;
        END
    END SE
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.231  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.250 6.865 2.630 ;
        RECT  6.525 2.010 6.865 2.630 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.689  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.250 0.790 13.590 4.140 ;
        RECT  11.810 2.190 13.590 2.630 ;
        RECT  11.810 0.790 12.150 4.140 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.970 -0.400 14.310 1.700 ;
        RECT  12.530 -0.400 12.870 1.700 ;
        RECT  11.090 -0.400 11.430 1.420 ;
        RECT  9.650 -0.400 9.990 1.495 ;
        RECT  8.210 -0.400 8.595 1.495 ;
        RECT  6.770 -0.400 7.110 1.495 ;
        RECT  5.090 -0.400 5.320 0.970 ;
        RECT  3.195 -0.400 3.480 1.320 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.970 2.720 14.310 5.280 ;
        RECT  12.530 3.290 12.870 5.280 ;
        RECT  11.090 2.940 11.430 5.280 ;
        RECT  8.790 2.940 9.130 5.280 ;
        RECT  5.845 3.520 6.830 5.280 ;
        RECT  2.730 2.670 3.380 3.010 ;
        RECT  2.730 2.670 3.030 5.280 ;
        RECT  0.740 2.720 1.045 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.505 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  1.275 2.120 1.505 4.210 ;
        RECT  1.275 3.870 2.040 4.210 ;
        RECT  0.180 0.830 0.520 1.170 ;
        RECT  0.180 0.940 2.345 1.170 ;
        RECT  1.735 0.940 2.345 1.280 ;
        RECT  1.735 0.940 1.965 3.065 ;
        RECT  1.735 2.725 2.230 3.065 ;
        RECT  4.170 1.090 4.400 2.350 ;
        RECT  2.870 2.010 4.550 2.350 ;
        RECT  4.210 2.010 4.550 3.010 ;
        RECT  3.710 0.630 4.860 0.860 ;
        RECT  5.550 0.630 6.185 0.950 ;
        RECT  4.630 0.630 4.860 1.430 ;
        RECT  5.550 0.630 5.780 1.430 ;
        RECT  4.630 1.200 5.780 1.430 ;
        RECT  3.710 0.630 3.940 1.780 ;
        RECT  2.195 1.550 3.940 1.780 ;
        RECT  2.195 1.510 2.535 1.850 ;
        RECT  4.865 1.200 5.095 3.780 ;
        RECT  4.865 3.440 5.425 3.780 ;
        RECT  6.010 1.310 6.295 2.010 ;
        RECT  5.325 1.660 6.295 2.010 ;
        RECT  5.845 1.660 6.185 2.970 ;
        RECT  8.930 1.155 9.270 2.490 ;
        RECT  10.370 1.155 10.710 2.490 ;
        RECT  7.490 1.155 7.830 2.370 ;
        RECT  7.640 2.150 11.580 2.490 ;
        RECT  7.640 2.150 7.980 3.860 ;
        RECT  9.940 2.150 10.280 3.860 ;
        RECT  0.180 0.940 1.30 1.170 ;
        RECT  7.640 2.150 10.70 2.490 ;
    END
END LSGCNX6

MACRO LSGCNX4
    CLASS CORE ;
    FOREIGN LSGCNX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.295 3.665 3.895 ;
        END
    END E
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 3.310 4.330 3.880 ;
        END
    END SE
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.550 1.840 7.440 2.180 ;
        RECT  6.425 2.250 6.805 2.630 ;
        RECT  6.550 1.840 6.805 2.630 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.017  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.420 2.250 11.790 2.630 ;
        RECT  11.450 0.780 11.790 2.630 ;
        RECT  10.730 2.250 11.070 3.880 ;
        RECT  9.420 2.240 10.350 2.630 ;
        RECT  10.010 1.230 10.350 2.630 ;
        RECT  9.210 2.970 9.720 3.880 ;
        RECT  9.420 2.240 9.720 3.880 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.730 -0.400 11.070 1.690 ;
        RECT  9.420 -0.400 9.760 0.710 ;
        RECT  8.100 -0.400 8.440 0.715 ;
        RECT  6.580 -0.400 6.920 0.710 ;
        RECT  5.100 -0.400 5.330 0.970 ;
        RECT  3.205 -0.400 3.490 1.320 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.450 2.970 11.790 5.280 ;
        RECT  9.970 2.970 10.310 5.280 ;
        RECT  8.490 2.970 8.830 5.280 ;
        RECT  5.485 3.540 6.360 5.280 ;
        RECT  2.730 2.670 3.380 3.010 ;
        RECT  2.730 2.670 3.030 5.280 ;
        RECT  0.740 2.720 1.045 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.505 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  1.275 2.120 1.505 4.210 ;
        RECT  1.275 3.870 2.040 4.210 ;
        RECT  0.180 0.830 0.520 1.170 ;
        RECT  0.180 0.940 2.350 1.170 ;
        RECT  1.735 0.940 2.350 1.280 ;
        RECT  1.735 0.940 1.965 3.065 ;
        RECT  1.735 2.725 2.230 3.065 ;
        RECT  4.180 1.090 4.410 2.350 ;
        RECT  2.870 2.010 4.550 2.350 ;
        RECT  4.210 2.010 4.550 3.010 ;
        RECT  3.720 0.630 4.870 0.860 ;
        RECT  5.560 0.630 6.185 0.970 ;
        RECT  4.640 0.630 4.870 1.430 ;
        RECT  5.560 0.630 5.790 1.430 ;
        RECT  4.640 1.200 5.790 1.430 ;
        RECT  3.720 0.630 3.950 1.780 ;
        RECT  2.195 1.550 3.950 1.780 ;
        RECT  2.195 1.510 2.535 1.850 ;
        RECT  4.780 1.200 5.065 3.810 ;
        RECT  4.725 3.470 5.065 3.810 ;
        RECT  6.020 1.330 6.320 2.000 ;
        RECT  5.325 1.660 6.320 2.000 ;
        RECT  5.325 1.660 5.765 2.990 ;
        RECT  7.340 1.150 9.000 1.490 ;
        RECT  8.660 1.150 9.000 2.710 ;
        RECT  8.660 2.370 9.190 2.710 ;
        RECT  7.340 2.410 9.190 2.710 ;
        RECT  7.340 2.410 7.680 3.880 ;
        RECT  0.180 0.940 1.10 1.170 ;
    END
END LSGCNX4

MACRO LSGCNX3
    CLASS CORE ;
    FOREIGN LSGCNX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.295 3.665 3.895 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.345  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.470 2.640 9.955 4.060 ;
        RECT  9.510 0.700 9.810 4.060 ;
        RECT  9.470 0.700 9.810 1.610 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 3.310 4.330 3.880 ;
        END
    END SE
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.698  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.030 7.710 2.630 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 1.610 ;
        RECT  8.750 -0.400 9.090 1.610 ;
        RECT  7.270 -0.400 7.630 0.960 ;
        RECT  5.240 -0.400 5.580 0.950 ;
        RECT  3.240 -0.400 3.525 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 2.640 10.530 5.280 ;
        RECT  8.750 2.640 9.090 5.280 ;
        RECT  6.570 3.440 6.910 5.280 ;
        RECT  5.470 3.480 5.810 5.280 ;
        RECT  2.730 2.670 3.380 3.010 ;
        RECT  2.730 2.670 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.485 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  1.255 2.120 1.485 4.210 ;
        RECT  1.255 3.870 1.825 4.210 ;
        RECT  0.180 0.830 0.520 1.170 ;
        RECT  1.715 0.765 2.350 1.105 ;
        RECT  0.180 0.940 1.945 1.170 ;
        RECT  1.715 0.765 1.945 3.065 ;
        RECT  1.715 2.725 2.230 3.065 ;
        RECT  2.870 1.795 4.550 2.210 ;
        RECT  4.215 1.090 4.550 3.010 ;
        RECT  4.210 1.795 4.550 3.010 ;
        RECT  3.755 0.630 5.010 0.860 ;
        RECT  6.040 0.630 6.380 0.970 ;
        RECT  4.780 0.630 5.010 3.780 ;
        RECT  6.040 0.630 6.295 1.410 ;
        RECT  4.780 1.180 6.295 1.410 ;
        RECT  3.755 0.630 3.985 1.565 ;
        RECT  2.175 1.335 3.985 1.565 ;
        RECT  2.175 1.335 2.500 1.840 ;
        RECT  4.780 1.180 5.050 3.780 ;
        RECT  4.710 3.440 5.050 3.780 ;
        RECT  6.525 1.270 7.010 1.610 ;
        RECT  6.525 1.270 6.825 1.930 ;
        RECT  6.030 1.640 6.825 1.930 ;
        RECT  6.030 1.640 6.370 3.040 ;
        RECT  8.030 1.880 9.280 2.220 ;
        RECT  8.030 0.700 8.370 4.240 ;
        RECT  7.760 3.900 8.370 4.240 ;
    END
END LSGCNX3

MACRO LSGCNX2
    CLASS CORE ;
    FOREIGN LSGCNX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.310 3.700 3.870 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.903  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.640 9.400 3.560 ;
        RECT  9.170 1.195 9.400 3.560 ;
        RECT  9.000 1.195 9.400 1.535 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.520  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 1.620 7.435 2.140 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.250 5.070 2.630 ;
        RECT  4.730 1.870 5.070 2.630 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  9.560 -0.400 9.900 0.710 ;
        RECT  8.280 -0.400 8.620 1.500 ;
        RECT  6.800 -0.400 7.160 0.930 ;
        RECT  5.205 -0.400 5.545 0.970 ;
        RECT  3.240 -0.400 3.525 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.560 3.960 9.900 5.280 ;
        RECT  8.280 2.640 8.620 5.280 ;
        RECT  5.510 3.475 5.850 5.280 ;
        RECT  2.730 2.615 3.380 2.955 ;
        RECT  2.730 2.615 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.485 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  1.255 2.120 1.485 4.210 ;
        RECT  1.255 3.870 1.825 4.210 ;
        RECT  0.180 0.830 0.520 1.170 ;
        RECT  1.715 0.765 2.350 1.105 ;
        RECT  0.180 0.940 1.945 1.170 ;
        RECT  1.715 0.765 1.945 3.065 ;
        RECT  1.715 2.725 2.230 3.065 ;
        RECT  4.215 1.090 4.515 1.430 ;
        RECT  4.215 1.090 4.500 2.020 ;
        RECT  2.870 1.795 4.305 2.210 ;
        RECT  4.050 1.795 4.305 3.780 ;
        RECT  4.050 3.440 4.390 3.780 ;
        RECT  3.755 0.630 4.975 0.860 ;
        RECT  5.775 0.630 6.420 0.970 ;
        RECT  4.745 0.630 4.975 1.430 ;
        RECT  4.745 1.200 6.005 1.430 ;
        RECT  3.755 0.630 3.985 1.565 ;
        RECT  2.175 1.335 3.985 1.565 ;
        RECT  2.175 1.335 2.500 1.840 ;
        RECT  5.775 0.630 6.005 3.245 ;
        RECT  4.750 2.905 6.005 3.245 ;
        RECT  6.235 1.280 6.690 4.100 ;
        RECT  7.560 1.040 7.905 1.380 ;
        RECT  7.665 1.880 8.860 2.220 ;
        RECT  7.665 1.040 7.905 2.900 ;
        RECT  7.130 2.560 7.905 2.900 ;
        RECT  7.130 2.560 7.470 3.880 ;
    END
END LSGCNX2

MACRO LSGCNX1
    CLASS CORE ;
    FOREIGN LSGCNX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.310 3.700 3.870 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.840 2.640 9.335 3.560 ;
        RECT  9.090 1.240 9.335 3.560 ;
        RECT  8.930 1.240 9.335 1.580 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.335  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.025 1.635 7.440 2.225 ;
        END
    END CLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.250 5.070 2.630 ;
        RECT  4.730 1.870 5.070 2.630 ;
        END
    END SE
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.360 -0.400 8.710 0.720 ;
        RECT  6.930 -0.400 7.275 1.050 ;
        RECT  5.205 -0.400 5.545 0.970 ;
        RECT  3.240 -0.400 3.525 0.970 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.130 2.920 8.460 5.280 ;
        RECT  5.710 3.650 6.050 5.280 ;
        RECT  2.730 2.615 3.380 2.955 ;
        RECT  2.730 2.615 3.030 5.280 ;
        RECT  0.740 2.720 1.025 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.400 0.520 2.460 ;
        RECT  0.180 2.120 1.485 2.460 ;
        RECT  0.180 1.400 0.510 3.800 ;
        RECT  1.255 2.120 1.485 4.210 ;
        RECT  1.255 3.870 1.825 4.210 ;
        RECT  0.180 0.830 0.520 1.170 ;
        RECT  1.715 0.765 2.350 1.105 ;
        RECT  0.180 0.940 1.945 1.170 ;
        RECT  1.715 0.765 1.945 3.065 ;
        RECT  1.715 2.725 2.230 3.065 ;
        RECT  4.215 1.090 4.515 1.430 ;
        RECT  4.215 1.090 4.500 2.020 ;
        RECT  2.870 1.795 4.305 2.210 ;
        RECT  4.050 1.795 4.305 3.780 ;
        RECT  4.050 3.440 4.390 3.780 ;
        RECT  3.755 0.630 4.975 0.860 ;
        RECT  5.775 0.630 6.420 0.970 ;
        RECT  4.745 0.630 4.975 1.430 ;
        RECT  4.745 1.200 6.005 1.430 ;
        RECT  3.755 0.630 3.985 1.565 ;
        RECT  2.175 1.335 3.985 1.565 ;
        RECT  2.175 1.335 2.500 1.840 ;
        RECT  5.775 0.630 6.005 3.245 ;
        RECT  4.950 2.905 6.005 3.245 ;
        RECT  6.235 1.310 6.670 3.210 ;
        RECT  7.670 0.710 8.020 2.220 ;
        RECT  7.670 1.880 8.860 2.220 ;
        RECT  7.670 0.710 7.900 3.170 ;
        RECT  6.970 2.830 7.900 3.170 ;
    END
END LSGCNX1

MACRO LSGCNX0
    CLASS CORE ;
    FOREIGN LSGCNX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.540 2.405 2.165 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.439  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.660 0.520 3.240 ;
        RECT  0.125 1.150 0.520 1.490 ;
        RECT  0.125 1.150 0.355 3.240 ;
        END
    END GCLK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.640 8.065 2.385 ;
        END
    END SE
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.100 6.995 2.630 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.320 -0.400 7.660 0.655 ;
        RECT  6.270 -0.400 6.610 0.655 ;
        RECT  4.810 -0.400 5.040 1.240 ;
        RECT  4.010 1.340 5.020 1.680 ;
        RECT  4.790 1.140 5.020 1.680 ;
        RECT  2.380 -0.400 3.260 0.870 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.300 4.035 8.640 5.280 ;
        RECT  6.380 3.720 6.720 5.280 ;
        RECT  3.940 3.550 4.280 5.280 ;
        RECT  3.010 3.720 3.350 5.280 ;
        RECT  0.980 2.660 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.555 1.025 1.920 1.310 ;
        RECT  1.555 1.025 1.900 1.340 ;
        RECT  0.630 1.815 0.970 2.155 ;
        RECT  0.630 1.925 1.785 2.155 ;
        RECT  1.555 1.025 1.785 2.980 ;
        RECT  1.555 2.640 2.550 2.980 ;
        RECT  2.940 1.270 3.295 1.610 ;
        RECT  2.940 1.270 3.225 3.480 ;
        RECT  2.210 3.250 3.225 3.480 ;
        RECT  2.210 3.250 2.550 3.780 ;
        RECT  3.525 0.630 4.580 0.940 ;
        RECT  3.485 1.760 3.755 1.930 ;
        RECT  3.525 0.630 3.755 1.930 ;
        RECT  3.455 1.785 3.685 3.175 ;
        RECT  3.455 2.880 5.225 3.175 ;
        RECT  4.890 2.880 5.225 3.365 ;
        RECT  4.890 2.880 5.175 3.370 ;
        RECT  3.915 2.100 5.245 2.440 ;
        RECT  5.935 1.345 7.455 1.635 ;
        RECT  5.935 1.345 6.220 1.955 ;
        RECT  7.225 1.345 7.455 3.220 ;
        RECT  7.225 2.880 8.010 3.220 ;
        RECT  7.890 0.630 8.360 0.865 ;
        RECT  7.890 0.630 8.125 1.115 ;
        RECT  5.475 0.885 8.125 1.115 ;
        RECT  5.250 1.340 5.705 1.680 ;
        RECT  5.330 3.570 5.705 3.905 ;
        RECT  5.475 0.885 5.705 3.905 ;
        RECT  5.325 3.620 5.705 3.905 ;
        RECT  8.355 1.095 8.705 1.435 ;
        RECT  7.500 3.575 8.705 3.805 ;
        RECT  8.475 1.095 8.705 3.805 ;
        RECT  6.955 3.775 7.840 4.115 ;
        RECT  5.475 0.885 7.30 1.115 ;
    END
END LSGCNX0

MACRO LOGIC1
    CLASS CORE ;
    FOREIGN LOGIC1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.629  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.430 1.135 3.250 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        RECT  0.180 3.780 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        RECT  0.400 -0.400 0.740 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.600 1.170 0.940 2.040 ;
        RECT  0.260 1.700 0.940 2.040 ;
    END
END LOGIC1

MACRO LOGIC0
    CLASS CORE ;
    FOREIGN LOGIC0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.418  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 1.030 1.135 1.690 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        RECT  0.400 3.650 0.740 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        RECT  0.180 -0.400 0.520 1.040 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.260 2.330 0.940 2.670 ;
        RECT  0.600 2.330 0.940 3.190 ;
    END
END LOGIC0

MACRO LGCPX8
    CLASS CORE ;
    FOREIGN LGCPX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.075 2.250 3.655 2.650 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.427  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.945 1.640 5.545 2.240 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.147  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.335 0.720 13.735 4.180 ;
        RECT  10.495 1.965 13.735 2.305 ;
        RECT  11.895 0.720 12.235 4.180 ;
        RECT  10.455 2.705 10.845 4.195 ;
        RECT  10.495 0.725 10.845 4.195 ;
        RECT  10.455 0.725 10.845 1.700 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.615 -0.400 12.955 1.700 ;
        RECT  11.175 -0.400 11.515 1.710 ;
        RECT  9.735 -0.400 10.080 1.555 ;
        RECT  7.435 -0.400 7.775 1.515 ;
        RECT  5.135 -0.400 5.475 1.410 ;
        RECT  3.150 -0.400 3.490 1.340 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.615 2.705 12.955 5.280 ;
        RECT  11.170 2.705 11.515 5.280 ;
        RECT  9.735 2.660 10.085 5.280 ;
        RECT  8.295 2.770 8.635 5.280 ;
        RECT  6.855 2.770 7.195 5.280 ;
        RECT  5.415 2.690 5.755 5.280 ;
        RECT  3.280 2.880 3.620 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 1.050 0.520 1.390 ;
        RECT  0.170 1.050 0.400 3.170 ;
        RECT  0.170 2.280 1.470 2.620 ;
        RECT  0.170 2.280 0.520 3.170 ;
        RECT  1.700 1.000 2.320 1.340 ;
        RECT  0.630 1.600 1.950 1.950 ;
        RECT  1.700 1.000 1.950 3.215 ;
        RECT  1.700 2.875 2.430 3.215 ;
        RECT  3.850 0.675 4.290 1.015 ;
        RECT  3.850 0.675 4.135 2.020 ;
        RECT  2.330 1.790 4.135 2.020 ;
        RECT  2.330 1.790 2.670 2.255 ;
        RECT  3.890 0.675 4.135 3.775 ;
        RECT  3.890 3.435 4.380 3.775 ;
        RECT  4.365 1.380 4.675 3.050 ;
        RECT  4.655 2.710 4.995 4.105 ;
        RECT  6.285 1.175 6.630 2.405 ;
        RECT  8.585 1.175 8.925 2.405 ;
        RECT  6.135 2.065 10.265 2.405 ;
        RECT  7.570 2.065 7.915 3.870 ;
        RECT  6.135 2.065 6.475 3.880 ;
        RECT  9.015 2.065 9.355 3.880 ;
        RECT  6.135 2.065 9.20 2.405 ;
    END
END LGCPX8

MACRO LGCPX6
    CLASS CORE ;
    FOREIGN LGCPX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.118  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.080 2.100 5.495 2.630 ;
        END
    END CLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.120 2.250 3.665 2.700 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.689  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.360 2.250 11.845 2.630 ;
        RECT  11.360 0.875 11.700 4.080 ;
        RECT  10.010 1.965 11.700 2.305 ;
        RECT  9.920 2.660 10.310 4.080 ;
        RECT  10.010 0.875 10.310 4.080 ;
        RECT  9.920 0.875 10.310 1.685 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.080 -0.400 12.420 1.630 ;
        RECT  10.640 -0.400 10.980 1.635 ;
        RECT  9.200 -0.400 9.545 1.555 ;
        RECT  6.855 -0.400 7.195 1.515 ;
        RECT  4.900 -0.400 5.245 0.900 ;
        RECT  3.380 -0.400 3.720 1.320 ;
        RECT  0.980 -0.400 1.320 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  12.080 2.660 12.420 5.280 ;
        RECT  10.635 2.660 10.980 5.280 ;
        RECT  9.200 2.660 9.525 5.280 ;
        RECT  7.760 2.770 8.100 5.280 ;
        RECT  6.320 2.745 6.660 5.280 ;
        RECT  4.840 3.480 5.180 5.280 ;
        RECT  3.320 3.480 3.610 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.240 1.470 2.580 ;
        RECT  0.180 0.980 0.520 3.170 ;
        RECT  1.630 1.000 2.520 1.345 ;
        RECT  1.630 1.000 1.930 1.920 ;
        RECT  0.750 1.570 1.930 1.920 ;
        RECT  1.700 1.000 1.930 3.215 ;
        RECT  1.700 2.875 2.430 3.215 ;
        RECT  3.950 0.890 4.525 1.230 ;
        RECT  3.950 0.890 4.180 1.910 ;
        RECT  2.330 1.680 4.180 1.910 ;
        RECT  2.330 1.680 2.890 2.210 ;
        RECT  2.660 1.680 2.890 3.250 ;
        RECT  2.660 3.020 4.045 3.250 ;
        RECT  3.840 3.110 4.070 3.820 ;
        RECT  3.840 3.480 4.380 3.820 ;
        RECT  4.900 1.360 5.240 1.700 ;
        RECT  4.465 1.460 5.240 1.700 ;
        RECT  4.090 2.140 4.695 2.480 ;
        RECT  4.465 1.460 4.695 3.000 ;
        RECT  4.275 2.140 4.695 3.000 ;
        RECT  5.705 1.270 6.045 1.555 ;
        RECT  5.725 1.270 6.045 2.405 ;
        RECT  8.030 1.175 8.370 2.405 ;
        RECT  5.725 2.065 9.780 2.405 ;
        RECT  5.725 1.270 5.955 3.330 ;
        RECT  5.600 2.995 5.955 3.330 ;
        RECT  8.475 2.065 8.820 3.545 ;
        RECT  7.040 2.065 7.380 3.555 ;
        RECT  5.725 2.065 8.80 2.405 ;
    END
END LGCPX6

MACRO LGCPX4
    CLASS CORE ;
    FOREIGN LGCPX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.120 2.250 3.665 2.700 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.515 1.640 6.175 2.185 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.254  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 1.200 10.585 3.910 ;
        RECT  8.840 1.965 10.585 2.305 ;
        RECT  8.750 2.660 9.140 3.910 ;
        RECT  8.840 1.200 9.140 3.910 ;
        RECT  8.750 1.200 9.140 1.540 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.545 ;
        RECT  8.030 -0.400 8.375 1.555 ;
        RECT  5.690 -0.400 6.030 1.340 ;
        RECT  4.890 -0.400 5.235 0.710 ;
        RECT  3.375 -0.400 3.715 1.340 ;
        RECT  0.980 -0.400 1.320 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.465 2.705 9.840 5.280 ;
        RECT  8.030 2.660 8.380 5.280 ;
        RECT  6.590 2.990 6.970 5.280 ;
        RECT  5.150 2.690 5.490 5.280 ;
        RECT  3.280 3.020 3.620 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.240 1.470 2.580 ;
        RECT  0.180 0.980 0.520 3.170 ;
        RECT  1.630 1.000 2.520 1.340 ;
        RECT  1.630 1.000 1.930 1.920 ;
        RECT  0.750 1.570 1.930 1.920 ;
        RECT  1.700 1.000 1.930 3.215 ;
        RECT  1.700 2.875 2.430 3.215 ;
        RECT  4.090 1.000 4.520 1.340 ;
        RECT  4.090 1.000 4.320 2.020 ;
        RECT  2.330 1.790 4.320 2.020 ;
        RECT  2.330 1.790 2.670 2.255 ;
        RECT  3.965 1.790 4.195 3.820 ;
        RECT  3.965 3.480 4.380 3.820 ;
        RECT  4.890 1.170 5.230 2.030 ;
        RECT  4.690 1.690 4.920 3.000 ;
        RECT  4.425 2.660 4.920 3.000 ;
        RECT  6.855 1.175 7.200 2.645 ;
        RECT  6.855 2.065 8.610 2.405 ;
        RECT  6.855 2.065 7.650 2.645 ;
        RECT  5.870 2.415 7.650 2.645 ;
        RECT  5.870 2.415 6.210 3.530 ;
        RECT  7.310 2.065 7.650 3.555 ;
    END
END LGCPX4

MACRO LGCPX3
    CLASS CORE ;
    FOREIGN LGCPX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.120 2.250 3.665 2.700 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.581  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.715 1.690 6.175 2.220 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.580 2.810 8.065 3.620 ;
        RECT  7.740 0.875 8.065 3.620 ;
        RECT  7.580 0.875 8.065 1.685 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.300 -0.400 8.640 1.635 ;
        RECT  6.865 -0.400 7.200 1.590 ;
        RECT  6.855 -0.400 7.200 1.105 ;
        RECT  4.890 -0.400 5.235 0.710 ;
        RECT  3.435 -0.400 3.775 1.340 ;
        RECT  0.980 -0.400 1.320 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.295 2.835 8.670 5.280 ;
        RECT  6.860 2.920 7.210 5.280 ;
        RECT  5.420 2.670 5.760 5.280 ;
        RECT  3.280 3.020 3.620 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.240 1.470 2.580 ;
        RECT  0.180 0.980 0.520 3.170 ;
        RECT  1.630 1.000 2.540 1.340 ;
        RECT  1.630 1.000 1.930 1.920 ;
        RECT  0.750 1.570 1.930 1.920 ;
        RECT  1.700 1.000 1.930 3.215 ;
        RECT  1.700 2.875 2.430 3.215 ;
        RECT  4.150 1.000 4.580 1.340 ;
        RECT  2.330 1.790 4.380 2.020 ;
        RECT  2.330 1.790 2.670 2.255 ;
        RECT  4.150 1.000 4.380 3.820 ;
        RECT  4.040 1.790 4.380 3.820 ;
        RECT  4.920 1.170 5.285 2.050 ;
        RECT  4.920 1.170 5.150 2.980 ;
        RECT  4.695 2.640 5.150 2.980 ;
        RECT  5.690 0.705 6.060 1.460 ;
        RECT  5.690 1.175 6.635 1.460 ;
        RECT  6.405 2.065 7.510 2.405 ;
        RECT  6.405 1.175 6.635 2.680 ;
        RECT  6.140 2.450 6.480 3.730 ;
        RECT  2.330 1.790 3.60 2.020 ;
    END
END LGCPX3

MACRO LGCPX2
    CLASS CORE ;
    FOREIGN LGCPX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.120 2.250 3.665 2.700 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.473  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.745 1.640 6.240 2.165 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.580 2.810 8.065 3.620 ;
        RECT  7.740 1.230 8.065 3.620 ;
        RECT  7.580 1.230 8.065 1.570 ;
        END
    END GCLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.300 -0.400 8.640 1.575 ;
        RECT  7.020 -0.400 7.360 0.710 ;
        RECT  4.945 -0.400 5.290 0.710 ;
        RECT  3.435 -0.400 3.775 1.340 ;
        RECT  0.980 -0.400 1.320 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.295 2.835 8.670 5.280 ;
        RECT  6.860 2.920 7.210 5.280 ;
        RECT  5.420 2.840 5.760 5.280 ;
        RECT  3.280 3.020 3.620 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.240 1.470 2.580 ;
        RECT  0.180 0.980 0.520 3.170 ;
        RECT  1.630 1.000 2.540 1.340 ;
        RECT  1.630 1.000 1.930 1.920 ;
        RECT  0.750 1.570 1.930 1.920 ;
        RECT  1.700 1.000 1.930 3.215 ;
        RECT  1.700 2.875 2.430 3.215 ;
        RECT  4.150 0.910 4.580 1.250 ;
        RECT  2.330 1.790 4.380 2.020 ;
        RECT  2.330 1.790 2.670 2.255 ;
        RECT  4.150 0.910 4.380 3.820 ;
        RECT  4.040 1.790 4.380 3.820 ;
        RECT  4.920 1.170 5.285 2.055 ;
        RECT  4.920 1.170 5.150 3.150 ;
        RECT  4.695 2.810 5.150 3.150 ;
        RECT  5.830 0.940 7.180 1.280 ;
        RECT  6.950 2.235 7.510 2.575 ;
        RECT  6.950 0.940 7.180 2.690 ;
        RECT  6.140 2.460 7.180 2.690 ;
        RECT  6.140 2.460 6.480 3.730 ;
        RECT  2.330 1.790 3.60 2.020 ;
    END
END LGCPX2

MACRO LGCPX1
    CLASS CORE ;
    FOREIGN LGCPX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.120 2.250 3.665 2.700 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 2.640 8.075 3.560 ;
        RECT  7.830 1.240 8.075 3.560 ;
        RECT  7.670 1.240 8.075 1.580 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.311  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.715 1.970 6.175 2.650 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.865 -0.400 7.215 1.555 ;
        RECT  4.945 -0.400 5.290 0.710 ;
        RECT  3.435 -0.400 3.775 1.340 ;
        RECT  0.980 -0.400 1.320 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.950 2.915 7.290 5.280 ;
        RECT  5.510 2.920 5.850 5.280 ;
        RECT  3.280 3.020 3.620 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.240 1.470 2.580 ;
        RECT  0.180 0.980 0.520 3.170 ;
        RECT  1.630 1.000 2.540 1.340 ;
        RECT  1.630 1.000 1.930 1.920 ;
        RECT  0.750 1.570 1.930 1.920 ;
        RECT  1.700 1.000 1.930 3.215 ;
        RECT  1.700 2.875 2.430 3.215 ;
        RECT  4.240 0.910 4.580 1.250 ;
        RECT  4.240 0.910 4.475 2.020 ;
        RECT  2.330 1.790 4.475 2.020 ;
        RECT  2.330 1.790 2.670 2.255 ;
        RECT  4.245 0.910 4.475 3.410 ;
        RECT  4.040 3.070 4.475 3.410 ;
        RECT  4.920 1.170 5.285 2.240 ;
        RECT  4.920 1.170 5.150 3.220 ;
        RECT  4.785 2.880 5.150 3.220 ;
        RECT  5.645 1.170 6.635 1.510 ;
        RECT  6.405 1.880 7.600 2.220 ;
        RECT  6.405 1.170 6.635 3.260 ;
        RECT  6.230 2.920 6.635 3.260 ;
        RECT  2.330 1.790 3.90 2.020 ;
    END
END LGCPX1

MACRO LGCPX0
    CLASS CORE ;
    FOREIGN LGCPX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.915 1.690 5.545 2.185 ;
        END
    END CLK
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.660 3.170 2.130 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 2.640 7.435 3.430 ;
        RECT  7.205 1.170 7.435 3.430 ;
        RECT  7.040 1.170 7.435 1.510 ;
        END
    END GCLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.240 2.640 6.580 5.280 ;
        RECT  4.765 3.750 5.105 5.280 ;
        RECT  4.790 3.725 5.105 5.280 ;
        RECT  3.085 2.900 3.425 5.280 ;
        RECT  0.980 2.780 1.320 5.280 ;
        RECT  0.610 2.780 1.320 3.120 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.240 -0.400 6.580 0.970 ;
        RECT  4.385 -0.400 4.725 0.710 ;
        RECT  2.870 -0.400 3.210 0.970 ;
        RECT  1.170 -0.400 1.455 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.195 1.105 0.480 2.360 ;
        RECT  0.195 2.070 1.230 2.360 ;
        RECT  0.135 2.125 0.365 4.060 ;
        RECT  0.135 3.720 0.520 4.060 ;
        RECT  0.475 0.630 0.940 0.875 ;
        RECT  1.700 0.630 2.165 0.970 ;
        RECT  0.710 0.630 0.940 1.785 ;
        RECT  0.710 1.555 1.930 1.785 ;
        RECT  1.700 0.630 1.930 3.120 ;
        RECT  1.700 2.830 2.180 3.120 ;
        RECT  3.655 0.630 4.035 0.970 ;
        RECT  2.160 1.200 3.885 1.430 ;
        RECT  2.160 1.200 2.415 2.470 ;
        RECT  3.655 0.630 3.885 3.055 ;
        RECT  3.655 2.715 4.225 3.055 ;
        RECT  4.385 1.170 4.725 1.510 ;
        RECT  4.385 1.170 4.685 2.030 ;
        RECT  4.115 1.690 4.685 2.030 ;
        RECT  4.455 1.170 4.685 3.520 ;
        RECT  3.965 3.290 4.685 3.520 ;
        RECT  3.965 3.290 4.305 3.760 ;
        RECT  5.210 1.170 6.005 1.460 ;
        RECT  6.590 1.815 6.930 2.155 ;
        RECT  5.775 1.925 6.930 2.155 ;
        RECT  5.775 1.170 6.005 3.180 ;
        RECT  5.435 2.840 6.005 3.180 ;
    END
END LGCPX0

MACRO LGCNX8
    CLASS CORE ;
    FOREIGN LGCNX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 1.640 3.655 2.020 ;
        RECT  2.960 1.640 3.300 2.210 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.857  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.455 2.035 13.735 2.335 ;
        RECT  13.335 0.700 13.735 2.335 ;
        RECT  12.615 2.035 12.955 3.770 ;
        RECT  11.895 0.700 12.235 2.335 ;
        RECT  11.295 2.035 11.635 3.770 ;
        RECT  9.975 2.745 10.795 3.085 ;
        RECT  10.455 1.130 10.795 3.085 ;
        RECT  9.975 2.745 10.315 3.770 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.633  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.800 6.025 2.140 ;
        RECT  5.165 1.800 5.545 2.630 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.615 -0.400 12.955 1.700 ;
        RECT  11.175 -0.400 11.515 1.805 ;
        RECT  9.895 -0.400 10.235 0.710 ;
        RECT  8.415 -0.400 8.755 1.280 ;
        RECT  6.975 -0.400 7.315 1.390 ;
        RECT  5.535 -0.400 5.875 1.390 ;
        RECT  3.240 -0.400 3.580 0.950 ;
        RECT  0.780 -0.400 1.120 0.740 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  13.335 2.735 13.675 5.280 ;
        RECT  12.055 4.170 12.395 5.280 ;
        RECT  10.735 4.170 11.075 5.280 ;
        RECT  9.415 4.170 9.755 5.280 ;
        RECT  7.075 2.840 7.415 5.280 ;
        RECT  4.070 3.540 5.075 5.280 ;
        RECT  2.460 2.530 3.380 2.870 ;
        RECT  2.460 2.530 2.800 5.280 ;
        RECT  0.740 2.645 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.060 0.520 2.350 ;
        RECT  0.180 2.010 1.320 2.350 ;
        RECT  0.180 1.060 0.510 4.060 ;
        RECT  1.630 0.630 2.350 0.950 ;
        RECT  1.630 0.630 1.930 2.980 ;
        RECT  1.630 2.640 2.230 2.980 ;
        RECT  1.485 2.700 1.825 4.150 ;
        RECT  3.885 0.630 4.380 0.970 ;
        RECT  2.175 1.180 4.115 1.410 ;
        RECT  2.175 1.180 2.515 1.840 ;
        RECT  3.885 0.630 4.115 2.480 ;
        RECT  3.610 2.250 4.115 2.480 ;
        RECT  3.610 2.250 3.840 3.780 ;
        RECT  3.085 3.440 3.840 3.780 ;
        RECT  4.740 0.630 5.080 1.570 ;
        RECT  4.345 1.200 5.080 1.570 ;
        RECT  4.345 1.200 4.675 3.050 ;
        RECT  4.175 2.710 4.675 3.050 ;
        RECT  7.695 0.940 8.035 2.610 ;
        RECT  9.135 0.940 9.475 2.490 ;
        RECT  6.255 1.050 6.595 2.610 ;
        RECT  6.255 2.270 10.225 2.490 ;
        RECT  7.695 2.150 10.225 2.490 ;
        RECT  5.925 2.370 8.565 2.610 ;
        RECT  5.925 2.370 6.265 3.880 ;
        RECT  8.225 2.150 8.565 3.880 ;
        RECT  6.255 2.270 9.80 2.490 ;
        RECT  7.695 2.150 9.20 2.490 ;
        RECT  5.925 2.370 7.80 2.610 ;
    END
END LGCNX8

MACRO LGCNX6
    CLASS CORE ;
    FOREIGN LGCNX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 1.640 3.655 2.020 ;
        RECT  2.960 1.640 3.300 2.210 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.974  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.615 2.035 13.105 2.630 ;
        RECT  12.615 2.035 12.955 3.770 ;
        RECT  10.455 2.035 13.105 2.335 ;
        RECT  11.895 0.700 12.235 2.335 ;
        RECT  11.295 2.035 11.635 3.770 ;
        RECT  9.975 2.745 10.795 3.085 ;
        RECT  10.455 1.130 10.795 3.085 ;
        RECT  9.975 2.745 10.315 3.770 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.238  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.800 6.025 2.140 ;
        RECT  5.165 1.800 5.545 2.630 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  12.615 -0.400 12.955 1.620 ;
        RECT  11.175 -0.400 11.515 1.620 ;
        RECT  9.895 -0.400 10.235 0.710 ;
        RECT  8.415 -0.400 8.755 1.280 ;
        RECT  6.975 -0.400 7.315 1.390 ;
        RECT  5.535 -0.400 5.875 1.390 ;
        RECT  3.240 -0.400 3.580 0.950 ;
        RECT  0.780 -0.400 1.120 0.740 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  12.055 4.170 12.395 5.280 ;
        RECT  10.735 4.170 11.075 5.280 ;
        RECT  9.415 4.170 9.755 5.280 ;
        RECT  7.075 3.000 7.415 5.280 ;
        RECT  4.070 3.540 5.075 5.280 ;
        RECT  2.460 2.530 3.380 2.870 ;
        RECT  2.460 2.530 2.800 5.280 ;
        RECT  0.740 2.645 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.060 0.520 2.350 ;
        RECT  0.180 2.010 1.320 2.350 ;
        RECT  0.180 1.060 0.510 4.060 ;
        RECT  1.630 0.630 2.350 0.950 ;
        RECT  1.630 0.630 1.930 2.980 ;
        RECT  1.630 2.640 2.230 2.980 ;
        RECT  1.485 2.700 1.825 4.150 ;
        RECT  3.885 0.630 4.380 0.970 ;
        RECT  2.175 1.180 4.115 1.410 ;
        RECT  2.175 1.180 2.515 1.840 ;
        RECT  3.885 0.630 4.115 2.480 ;
        RECT  3.610 2.250 4.115 2.480 ;
        RECT  3.610 2.250 3.840 3.780 ;
        RECT  3.085 3.440 3.840 3.780 ;
        RECT  4.740 0.630 5.080 1.570 ;
        RECT  4.345 1.200 5.080 1.570 ;
        RECT  4.345 1.200 4.675 3.050 ;
        RECT  4.175 2.710 4.675 3.050 ;
        RECT  7.695 0.940 8.035 2.610 ;
        RECT  9.135 0.940 9.475 2.490 ;
        RECT  6.255 1.050 6.595 2.610 ;
        RECT  6.255 2.270 10.225 2.490 ;
        RECT  7.695 2.150 10.225 2.490 ;
        RECT  5.925 2.370 8.565 2.610 ;
        RECT  5.925 2.370 6.265 3.880 ;
        RECT  8.225 2.150 8.565 3.880 ;
        RECT  6.255 2.270 9.30 2.490 ;
        RECT  7.695 2.150 9.70 2.490 ;
        RECT  5.925 2.370 7.30 2.610 ;
    END
END LGCNX6

MACRO LGCNX4
    CLASS CORE ;
    FOREIGN LGCNX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 1.640 3.655 2.020 ;
        RECT  2.960 1.640 3.300 2.210 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.046  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.160 2.250 10.530 2.630 ;
        RECT  10.190 0.710 10.530 2.630 ;
        RECT  9.470 2.250 9.810 3.780 ;
        RECT  8.750 1.320 9.090 2.630 ;
        RECT  7.950 2.910 8.460 3.780 ;
        RECT  8.160 2.250 8.460 3.780 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.850 6.180 2.190 ;
        RECT  5.165 1.850 5.545 2.630 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.700 ;
        RECT  8.160 -0.400 8.500 0.880 ;
        RECT  6.840 -0.400 7.180 0.715 ;
        RECT  5.520 -0.400 5.860 0.710 ;
        RECT  3.240 -0.400 3.580 0.950 ;
        RECT  0.780 -0.400 1.120 0.740 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 2.860 10.530 5.280 ;
        RECT  8.710 2.860 9.050 5.280 ;
        RECT  7.230 2.910 7.570 5.280 ;
        RECT  4.070 3.540 5.270 5.280 ;
        RECT  2.460 2.530 3.380 2.870 ;
        RECT  2.460 2.530 2.800 5.280 ;
        RECT  0.740 2.645 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.060 0.520 2.350 ;
        RECT  0.180 2.010 1.320 2.350 ;
        RECT  0.180 1.060 0.510 4.060 ;
        RECT  1.630 0.630 2.350 0.950 ;
        RECT  1.630 0.630 1.930 2.980 ;
        RECT  1.630 2.640 2.230 2.980 ;
        RECT  1.485 2.700 1.825 4.150 ;
        RECT  3.885 0.630 4.380 0.970 ;
        RECT  2.175 1.180 4.115 1.410 ;
        RECT  2.175 1.180 2.515 1.840 ;
        RECT  3.885 0.630 4.115 2.480 ;
        RECT  3.610 2.250 4.115 2.480 ;
        RECT  3.610 2.250 3.840 3.780 ;
        RECT  3.085 3.440 3.840 3.780 ;
        RECT  4.820 0.630 5.160 1.500 ;
        RECT  4.345 1.200 5.160 1.500 ;
        RECT  4.345 1.200 4.690 1.550 ;
        RECT  4.345 1.200 4.675 2.970 ;
        RECT  4.330 2.630 4.675 2.970 ;
        RECT  6.080 1.280 6.640 1.620 ;
        RECT  6.410 1.280 6.640 2.660 ;
        RECT  7.400 1.280 7.740 2.660 ;
        RECT  6.410 2.270 7.930 2.660 ;
        RECT  6.080 2.420 6.420 3.880 ;
    END
END LGCNX4

MACRO LGCNX3
    CLASS CORE ;
    FOREIGN LGCNX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 1.640 3.655 2.020 ;
        RECT  2.960 1.640 3.300 2.210 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.560  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 2.840 9.270 3.760 ;
        RECT  7.610 2.840 9.270 3.240 ;
        RECT  7.855 0.700 8.195 3.240 ;
        RECT  7.610 2.840 7.950 3.760 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.689  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.930 5.545 2.630 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.575 -0.400 8.915 1.620 ;
        RECT  7.135 -0.400 7.475 1.620 ;
        RECT  5.695 -0.400 6.040 1.620 ;
        RECT  3.240 -0.400 3.580 0.950 ;
        RECT  0.780 -0.400 1.120 0.740 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.050 4.160 8.510 5.280 ;
        RECT  4.070 3.480 5.010 5.280 ;
        RECT  2.460 2.530 3.380 2.870 ;
        RECT  2.460 2.530 2.800 5.280 ;
        RECT  0.740 2.645 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.060 0.520 2.350 ;
        RECT  0.180 2.010 1.320 2.350 ;
        RECT  0.180 1.060 0.510 4.060 ;
        RECT  1.630 0.630 2.350 0.950 ;
        RECT  1.630 0.630 1.930 2.980 ;
        RECT  1.630 2.640 2.230 2.980 ;
        RECT  1.485 2.700 1.825 4.150 ;
        RECT  3.885 0.630 4.380 0.970 ;
        RECT  2.175 1.180 4.115 1.410 ;
        RECT  2.175 1.180 2.515 1.840 ;
        RECT  3.885 0.630 4.115 2.480 ;
        RECT  3.610 2.250 4.115 2.480 ;
        RECT  3.610 2.250 3.840 3.780 ;
        RECT  3.085 3.440 3.840 3.780 ;
        RECT  4.345 1.280 5.235 1.620 ;
        RECT  4.345 1.280 4.675 3.040 ;
        RECT  4.110 2.710 4.675 3.040 ;
        RECT  6.415 0.700 6.755 2.610 ;
        RECT  5.860 2.270 7.625 2.610 ;
        RECT  5.860 2.270 6.200 3.760 ;
    END
END LGCNX3

MACRO LGCNX2
    CLASS CORE ;
    FOREIGN LGCNX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.300 2.210 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.906  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 2.640 7.450 3.560 ;
        RECT  7.220 1.160 7.450 3.560 ;
        RECT  7.110 1.160 7.450 1.500 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.520  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.010 1.640 5.545 2.110 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 0.710 ;
        RECT  6.390 -0.400 6.730 1.470 ;
        RECT  4.910 -0.400 5.255 0.940 ;
        RECT  3.240 -0.400 3.580 0.950 ;
        RECT  0.780 -0.400 1.120 0.740 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.680 2.640 8.010 5.280 ;
        RECT  6.230 2.645 6.570 5.280 ;
        RECT  3.820 3.910 4.160 5.280 ;
        RECT  2.460 2.480 3.380 2.820 ;
        RECT  2.460 2.480 2.800 5.280 ;
        RECT  0.740 2.720 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.060 0.520 2.350 ;
        RECT  0.180 2.010 1.270 2.350 ;
        RECT  0.180 1.060 0.510 4.060 ;
        RECT  1.545 0.630 2.350 0.950 ;
        RECT  1.545 0.630 1.845 4.150 ;
        RECT  1.545 2.640 2.230 2.980 ;
        RECT  1.545 2.640 1.885 4.150 ;
        RECT  3.810 0.630 4.380 0.970 ;
        RECT  3.810 0.630 4.040 1.410 ;
        RECT  2.075 1.180 4.040 1.410 ;
        RECT  2.075 1.180 2.415 1.840 ;
        RECT  3.610 1.180 3.840 3.680 ;
        RECT  3.060 3.440 3.840 3.680 ;
        RECT  3.060 3.440 3.400 3.780 ;
        RECT  4.270 1.340 4.720 2.460 ;
        RECT  4.070 2.120 4.720 2.460 ;
        RECT  4.380 1.340 4.720 3.470 ;
        RECT  5.670 1.070 6.130 1.410 ;
        RECT  5.775 1.070 6.130 2.210 ;
        RECT  5.775 1.870 6.990 2.210 ;
        RECT  5.775 1.070 6.005 2.595 ;
        RECT  5.080 2.365 6.005 2.595 ;
        RECT  5.080 2.365 5.420 3.880 ;
    END
END LGCNX2

MACRO LGCNX1
    CLASS CORE ;
    FOREIGN LGCNX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 1.640 3.655 2.210 ;
        END
    END E
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 2.640 7.445 3.560 ;
        RECT  7.200 1.270 7.445 3.560 ;
        RECT  7.040 1.270 7.445 1.610 ;
        END
    END GCLK
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.335  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.135 1.635 5.550 2.220 ;
        END
    END CLK
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.470 -0.400 6.820 0.720 ;
        RECT  5.040 -0.400 5.385 1.050 ;
        RECT  3.240 -0.400 3.580 0.950 ;
        RECT  0.780 -0.400 1.120 0.740 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.230 2.780 6.570 5.280 ;
        RECT  3.820 3.910 4.160 5.280 ;
        RECT  2.460 2.480 3.380 2.820 ;
        RECT  2.460 2.480 2.800 5.280 ;
        RECT  0.740 2.720 1.080 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.060 0.520 2.350 ;
        RECT  0.180 2.010 1.320 2.350 ;
        RECT  0.180 1.060 0.510 4.060 ;
        RECT  1.630 0.630 2.350 0.950 ;
        RECT  1.630 0.630 1.930 2.980 ;
        RECT  1.630 2.640 2.230 2.980 ;
        RECT  1.485 2.700 1.825 4.150 ;
        RECT  3.885 0.630 4.380 0.970 ;
        RECT  2.160 1.180 4.115 1.410 ;
        RECT  2.160 1.180 2.500 1.840 ;
        RECT  3.885 0.630 4.115 3.680 ;
        RECT  3.060 3.440 4.115 3.680 ;
        RECT  3.060 3.440 3.400 3.780 ;
        RECT  4.345 1.310 4.780 3.470 ;
        RECT  5.780 0.710 6.130 2.220 ;
        RECT  5.780 1.880 6.970 2.220 ;
        RECT  5.780 0.710 6.010 2.680 ;
        RECT  5.080 2.450 6.010 2.680 ;
        RECT  5.080 2.450 5.420 3.170 ;
    END
END LGCNX1

MACRO LGCNX0
    CLASS CORE ;
    FOREIGN LGCNX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.660 3.125 2.255 ;
        END
    END E
    PIN CLK
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 3.300 6.175 3.850 ;
        RECT  5.345 3.300 6.175 3.640 ;
        RECT  5.300 3.300 6.175 3.625 ;
        END
    END CLK
    PIN GCLK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 2.285 7.435 2.980 ;
        RECT  7.160 1.170 7.435 2.980 ;
        RECT  7.040 1.170 7.435 1.510 ;
        END
    END GCLK
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.405 2.640 6.745 5.280 ;
        RECT  6.240 2.640 6.745 2.980 ;
        RECT  4.765 3.750 5.105 5.280 ;
        RECT  4.785 3.720 5.090 5.280 ;
        RECT  3.070 2.840 3.410 5.280 ;
        RECT  1.075 2.720 1.415 5.280 ;
        RECT  0.595 2.720 1.415 3.060 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.240 -0.400 6.580 0.870 ;
        RECT  5.040 -0.400 5.380 0.870 ;
        RECT  2.855 -0.400 3.195 0.970 ;
        RECT  0.795 -0.400 1.135 0.760 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.135 1.060 0.535 1.400 ;
        RECT  0.135 2.010 1.215 2.300 ;
        RECT  0.135 1.060 0.365 4.030 ;
        RECT  0.135 3.690 0.845 4.030 ;
        RECT  1.645 1.270 1.930 3.750 ;
        RECT  1.645 2.720 2.165 3.060 ;
        RECT  1.645 2.720 1.985 3.750 ;
        RECT  3.640 0.630 4.020 0.915 ;
        RECT  2.160 1.200 3.870 1.430 ;
        RECT  2.160 1.200 2.415 2.100 ;
        RECT  3.640 0.630 3.870 3.055 ;
        RECT  3.640 2.715 4.210 3.055 ;
        RECT  4.230 1.245 4.570 2.110 ;
        RECT  4.100 1.770 4.670 2.110 ;
        RECT  4.440 1.770 4.670 3.520 ;
        RECT  3.965 3.290 4.670 3.520 ;
        RECT  3.965 3.290 4.305 3.760 ;
        RECT  5.640 1.170 6.005 1.510 ;
        RECT  5.775 1.740 6.930 2.055 ;
        RECT  5.775 1.170 6.005 3.055 ;
        RECT  5.010 2.715 6.005 3.055 ;
    END
END LGCNX0

MACRO ITLX8
    CLASS CORE ;
    FOREIGN ITLX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.720  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.930 2.250 6.805 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 5.573  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.075 0.700 12.475 4.180 ;
        RECT  7.750 1.870 12.475 2.370 ;
        RECT  12.070 0.700 12.475 2.370 ;
        RECT  10.635 0.700 10.980 2.370 ;
        RECT  10.635 0.700 10.975 4.180 ;
        RECT  9.195 0.700 9.545 2.370 ;
        RECT  9.195 0.700 9.535 4.180 ;
        RECT  7.750 0.700 8.090 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.716  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.710 4.190 ;
        END
    END EN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.360 -0.400 11.700 1.600 ;
        RECT  9.920 -0.400 10.260 1.600 ;
        RECT  8.475 -0.400 8.815 1.600 ;
        RECT  6.950 -0.400 7.290 0.940 ;
        RECT  5.245 -0.400 5.585 1.020 ;
        RECT  3.805 -0.400 4.145 1.075 ;
        RECT  0.945 -0.400 1.285 1.620 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.355 2.640 11.695 5.280 ;
        RECT  9.915 2.640 10.255 5.280 ;
        RECT  8.470 2.640 8.810 5.280 ;
        RECT  6.935 3.840 7.275 5.280 ;
        RECT  5.335 3.840 5.700 5.280 ;
        RECT  3.900 3.320 4.240 5.280 ;
        RECT  0.940 2.800 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.230 1.430 2.570 ;
        RECT  0.180 1.175 0.520 3.220 ;
        RECT  6.105 1.635 6.445 1.970 ;
        RECT  5.345 1.740 6.445 1.970 ;
        RECT  5.345 1.740 5.580 2.410 ;
        RECT  4.320 2.070 5.580 2.410 ;
        RECT  5.350 1.740 5.580 3.150 ;
        RECT  5.350 2.865 6.450 3.150 ;
        RECT  2.385 1.150 2.725 1.995 ;
        RECT  2.385 1.765 3.520 1.995 ;
        RECT  3.180 2.860 4.980 3.090 ;
        RECT  4.620 2.860 4.980 3.610 ;
        RECT  7.190 2.310 7.520 3.610 ;
        RECT  4.620 3.380 7.520 3.610 ;
        RECT  1.660 2.755 2.000 4.250 ;
        RECT  4.620 2.860 4.960 4.185 ;
        RECT  3.180 1.765 3.520 4.250 ;
        RECT  1.660 4.020 3.520 4.250 ;
        RECT  1.665 0.630 3.425 0.885 ;
        RECT  4.525 0.700 4.865 1.650 ;
        RECT  3.085 0.630 3.425 1.535 ;
        RECT  4.525 1.250 7.520 1.405 ;
        RECT  5.760 1.170 7.520 1.405 ;
        RECT  3.085 1.305 5.930 1.480 ;
        RECT  3.085 1.305 4.870 1.535 ;
        RECT  4.525 1.250 4.870 1.650 ;
        RECT  7.225 1.170 7.520 1.980 ;
        RECT  1.665 0.630 2.005 2.455 ;
        RECT  1.665 2.225 2.720 2.455 ;
        RECT  2.380 2.225 2.720 3.790 ;
        RECT  4.620 3.380 6.70 3.610 ;
        RECT  4.525 1.250 6.90 1.405 ;
        RECT  3.085 1.305 4.70 1.480 ;
    END
END ITLX8

MACRO ITLX6
    CLASS CORE ;
    FOREIGN ITLX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.055 6.325 2.340 ;
        RECT  5.795 2.055 6.210 2.580 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.180 0.700 10.585 4.180 ;
        RECT  7.300 1.870 10.585 2.210 ;
        RECT  10.175 0.700 10.585 2.210 ;
        RECT  8.740 0.700 9.085 2.210 ;
        RECT  8.740 0.700 9.080 4.180 ;
        RECT  7.300 0.700 7.650 2.210 ;
        RECT  7.300 0.700 7.640 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.460 2.595 2.230 2.940 ;
        RECT  1.460 1.610 1.690 2.940 ;
        RECT  0.755 1.610 1.690 2.020 ;
        END
    END EN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.460 2.740 9.800 5.280 ;
        RECT  8.020 2.740 8.360 5.280 ;
        RECT  6.580 2.730 6.920 5.280 ;
        RECT  5.120 3.270 5.460 5.280 ;
        RECT  3.680 3.255 4.020 5.280 ;
        RECT  0.760 4.070 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.465 -0.400 9.805 1.575 ;
        RECT  8.025 -0.400 8.365 1.570 ;
        RECT  6.580 -0.400 6.920 1.365 ;
        RECT  3.825 -0.400 5.125 0.975 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.280 1.230 2.620 ;
        RECT  0.180 1.090 0.520 3.570 ;
        RECT  2.380 1.360 2.720 1.905 ;
        RECT  2.380 1.675 3.150 1.905 ;
        RECT  2.920 1.675 3.150 4.130 ;
        RECT  2.920 2.660 3.335 3.025 ;
        RECT  2.920 2.795 4.740 3.025 ;
        RECT  1.520 3.195 1.860 4.130 ;
        RECT  4.400 2.795 4.740 3.880 ;
        RECT  2.920 2.660 3.300 4.130 ;
        RECT  1.520 3.790 3.300 4.130 ;
        RECT  4.155 2.205 5.525 2.545 ;
        RECT  5.275 2.205 5.525 3.040 ;
        RECT  5.275 2.810 6.160 3.040 ;
        RECT  5.820 2.810 6.160 3.880 ;
        RECT  5.330 1.080 6.205 1.365 ;
        RECT  1.620 0.900 3.595 1.130 ;
        RECT  1.620 0.900 2.150 1.240 ;
        RECT  3.365 0.900 3.595 1.580 ;
        RECT  3.380 1.350 5.100 1.695 ;
        RECT  4.850 1.595 7.070 1.825 ;
        RECT  6.760 1.595 7.070 2.100 ;
        RECT  1.920 0.900 2.150 2.365 ;
        RECT  1.920 2.135 2.690 2.365 ;
        RECT  2.460 2.135 2.690 3.515 ;
        RECT  2.240 3.170 2.690 3.515 ;
        RECT  4.850 1.595 6.80 1.825 ;
    END
END ITLX6

MACRO ITLX4
    CLASS CORE ;
    FOREIGN ITLX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.356  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.795 2.165 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.575 0.995 8.065 4.120 ;
        RECT  6.135 1.840 8.065 2.175 ;
        RECT  6.135 0.995 6.485 2.175 ;
        RECT  6.135 0.995 6.475 4.120 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 2.640 2.050 2.985 ;
        RECT  1.415 1.545 1.645 2.985 ;
        RECT  0.755 1.545 1.645 1.990 ;
        END
    END EN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.295 2.800 8.635 5.280 ;
        RECT  6.855 2.800 7.195 5.280 ;
        RECT  5.415 2.800 5.755 5.280 ;
        RECT  3.935 2.855 5.755 3.085 ;
        RECT  3.935 2.855 4.275 3.790 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.300 -0.400 8.640 1.335 ;
        RECT  6.860 -0.400 7.200 1.335 ;
        RECT  5.415 -0.400 5.755 1.435 ;
        RECT  3.900 -0.400 4.240 0.950 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.220 1.185 2.560 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.540 0.785 2.960 1.125 ;
        RECT  1.885 0.785 2.960 1.130 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.570 2.410 ;
        RECT  2.280 2.180 2.570 3.515 ;
        RECT  3.190 1.050 3.480 1.410 ;
        RECT  3.190 1.180 4.255 1.410 ;
        RECT  4.025 1.880 4.515 2.220 ;
        RECT  4.025 1.180 4.255 2.625 ;
        RECT  3.260 2.395 4.255 2.625 ;
        RECT  3.260 2.395 3.555 3.790 ;
        RECT  2.345 1.360 2.640 1.950 ;
        RECT  2.345 1.720 3.030 1.950 ;
        RECT  1.520 3.245 1.860 4.085 ;
        RECT  2.800 1.720 3.030 4.250 ;
        RECT  1.520 3.745 3.030 4.085 ;
        RECT  4.655 3.315 4.995 4.250 ;
        RECT  2.800 4.020 4.995 4.250 ;
        RECT  4.660 1.105 5.000 1.450 ;
        RECT  4.750 1.105 5.000 2.110 ;
        RECT  4.750 1.880 5.905 2.110 ;
        RECT  5.570 1.880 5.905 2.220 ;
        RECT  2.800 4.020 3.30 4.250 ;
    END
END ITLX4

MACRO ITLX3
    CLASS CORE ;
    FOREIGN ITLX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.425 2.640 2.050 2.985 ;
        RECT  1.425 1.765 1.655 2.985 ;
        RECT  0.755 1.765 1.655 1.995 ;
        RECT  0.755 1.545 1.230 1.995 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.460 3.755 4.085 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.625 2.250 8.065 2.630 ;
        RECT  7.625 0.995 7.970 3.965 ;
        RECT  6.185 1.840 7.970 2.180 ;
        RECT  6.185 0.995 6.535 2.180 ;
        RECT  6.185 0.995 6.525 3.965 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.905 2.645 7.245 5.280 ;
        RECT  5.425 2.520 5.805 5.280 ;
        RECT  3.985 2.520 4.325 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.910 -0.400 7.250 1.335 ;
        RECT  5.465 -0.400 5.805 1.335 ;
        RECT  3.985 -0.400 4.325 1.390 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.225 1.195 2.565 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.880 0.785 3.040 1.130 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.585 2.410 ;
        RECT  2.280 2.180 2.585 3.255 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.045 1.950 ;
        RECT  1.520 3.245 1.860 3.825 ;
        RECT  2.815 1.720 3.045 3.825 ;
        RECT  1.520 3.485 3.045 3.825 ;
        RECT  3.275 1.870 4.565 2.210 ;
        RECT  3.275 1.020 3.605 3.125 ;
        RECT  4.705 2.520 5.045 4.250 ;
        RECT  4.705 1.105 5.045 1.450 ;
        RECT  4.795 1.105 5.045 2.040 ;
        RECT  4.795 1.700 5.955 2.040 ;
    END
END ITLX3

MACRO ITLX20
    CLASS CORE ;
    FOREIGN ITLX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.720 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.667  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.285 2.070 14.030 2.410 ;
        RECT  13.350 2.070 13.745 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  27.200 0.700 27.595 4.180 ;
        RECT  16.810 1.840 27.595 2.490 ;
        RECT  25.760 0.700 26.100 4.180 ;
        RECT  25.750 0.700 26.100 2.490 ;
        RECT  24.320 0.700 24.665 4.180 ;
        RECT  24.310 0.700 24.665 2.490 ;
        RECT  22.880 0.700 23.220 4.180 ;
        RECT  22.875 0.700 23.220 2.490 ;
        RECT  21.440 0.700 21.780 4.180 ;
        RECT  21.435 0.700 21.780 2.490 ;
        RECT  20.000 0.700 20.350 2.490 ;
        RECT  20.000 0.700 20.340 4.180 ;
        RECT  18.560 0.700 18.900 4.180 ;
        RECT  17.120 0.700 17.460 4.180 ;
        RECT  15.680 2.810 17.460 3.090 ;
        RECT  16.810 1.155 17.460 3.090 ;
        RECT  15.600 1.155 17.460 1.385 ;
        RECT  15.680 2.810 16.020 4.180 ;
        RECT  15.600 0.850 15.940 1.385 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.768  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.880 0.530 2.630 ;
        END
    END EN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 27.720 0.400 ;
        RECT  26.480 -0.400 26.820 1.570 ;
        RECT  25.040 -0.400 25.380 1.570 ;
        RECT  23.600 -0.400 23.940 1.575 ;
        RECT  22.160 -0.400 22.500 1.570 ;
        RECT  20.720 -0.400 21.060 1.570 ;
        RECT  19.280 -0.400 19.620 1.570 ;
        RECT  17.840 -0.400 18.180 1.570 ;
        RECT  16.355 -0.400 16.700 0.925 ;
        RECT  14.765 -0.400 15.105 1.195 ;
        RECT  11.520 -0.400 13.245 0.655 ;
        RECT  10.260 -0.400 10.600 1.510 ;
        RECT  8.820 -0.400 9.160 1.510 ;
        RECT  7.380 -0.400 7.720 1.140 ;
        RECT  5.940 -0.400 6.280 1.075 ;
        RECT  3.060 -0.400 3.400 1.285 ;
        RECT  1.620 -0.400 1.960 1.385 ;
        RECT  0.180 -0.400 0.520 1.650 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 27.720 5.280 ;
        RECT  26.480 2.760 26.820 5.280 ;
        RECT  25.040 2.760 25.380 5.280 ;
        RECT  23.600 2.760 23.940 5.280 ;
        RECT  22.160 2.760 22.500 5.280 ;
        RECT  20.720 2.760 21.060 5.280 ;
        RECT  19.280 2.760 19.620 5.280 ;
        RECT  17.840 2.760 18.180 5.280 ;
        RECT  16.400 3.320 16.740 5.280 ;
        RECT  14.440 3.840 15.300 5.280 ;
        RECT  14.960 2.810 15.300 5.280 ;
        RECT  12.960 3.840 13.300 5.280 ;
        RECT  11.520 3.840 11.860 5.280 ;
        RECT  10.260 3.200 10.600 5.280 ;
        RECT  8.820 3.200 9.160 5.280 ;
        RECT  7.380 3.200 7.720 5.280 ;
        RECT  5.940 3.200 6.280 5.280 ;
        RECT  3.060 3.220 3.400 5.280 ;
        RECT  1.620 2.765 1.960 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.140 2.440 2.480 ;
        RECT  0.900 0.830 1.240 3.910 ;
        RECT  11.755 1.345 14.005 1.655 ;
        RECT  5.705 2.070 7.960 2.460 ;
        RECT  5.705 2.200 12.055 2.460 ;
        RECT  11.755 1.345 12.055 3.150 ;
        RECT  11.755 2.830 12.580 3.150 ;
        RECT  11.755 2.860 14.030 3.150 ;
        RECT  4.500 1.115 4.840 1.995 ;
        RECT  4.500 1.765 5.450 1.995 ;
        RECT  14.260 2.230 16.380 2.570 ;
        RECT  5.220 1.765 5.450 4.250 ;
        RECT  5.220 2.690 11.320 2.970 ;
        RECT  2.340 2.710 4.120 2.990 ;
        RECT  10.980 2.690 11.320 3.610 ;
        RECT  14.260 2.230 14.560 3.610 ;
        RECT  10.980 3.380 14.560 3.610 ;
        RECT  2.340 2.710 2.680 3.680 ;
        RECT  3.780 2.710 4.120 4.250 ;
        RECT  6.660 2.690 7.000 4.120 ;
        RECT  8.100 2.690 8.445 4.120 ;
        RECT  9.540 2.690 9.880 4.145 ;
        RECT  5.220 2.690 5.560 4.250 ;
        RECT  3.780 3.970 5.560 4.250 ;
        RECT  3.780 0.630 5.560 0.885 ;
        RECT  10.980 0.885 14.535 1.115 ;
        RECT  5.220 0.630 5.560 1.535 ;
        RECT  6.660 0.730 7.000 1.650 ;
        RECT  2.340 0.945 2.680 1.795 ;
        RECT  5.220 1.305 7.000 1.535 ;
        RECT  14.260 0.885 14.535 1.900 ;
        RECT  8.100 0.740 8.440 1.650 ;
        RECT  6.660 1.370 8.440 1.650 ;
        RECT  8.170 0.740 8.440 1.970 ;
        RECT  9.540 0.740 9.880 1.970 ;
        RECT  3.780 0.630 4.120 1.795 ;
        RECT  2.340 1.515 4.120 1.795 ;
        RECT  14.260 1.615 16.385 1.900 ;
        RECT  10.980 0.885 11.320 1.970 ;
        RECT  8.170 1.740 11.320 1.970 ;
        RECT  3.790 0.630 4.120 2.455 ;
        RECT  3.790 2.225 4.840 2.455 ;
        RECT  4.500 2.225 4.840 3.740 ;
        RECT  11.755 1.345 13.20 1.655 ;
        RECT  5.705 2.070 6.80 2.460 ;
        RECT  5.705 2.200 11.60 2.460 ;
        RECT  11.755 2.860 13.40 3.150 ;
        RECT  14.260 2.230 15.90 2.570 ;
        RECT  5.220 2.690 10.40 2.970 ;
        RECT  10.980 3.380 13.60 3.610 ;
        RECT  10.980 0.885 13.50 1.115 ;
        RECT  14.260 1.615 15.30 1.900 ;
        RECT  8.170 1.740 10.40 1.970 ;
    END
END ITLX20

MACRO ITLX2
    CLASS CORE ;
    FOREIGN ITLX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.460 3.760 4.085 ;
        END
    END A
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.425 2.640 2.110 2.985 ;
        RECT  1.425 1.545 1.655 2.985 ;
        RECT  0.755 1.545 1.655 2.020 ;
        END
    END EN
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.084  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.945 0.995 7.435 3.965 ;
        RECT  5.505 1.840 7.435 2.180 ;
        RECT  5.505 0.995 5.855 2.180 ;
        RECT  5.505 0.995 5.845 3.680 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.225 2.645 6.565 5.280 ;
        RECT  4.025 2.640 4.365 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.230 -0.400 6.570 1.335 ;
        RECT  4.025 -0.400 4.365 1.585 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.250 1.195 2.555 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.880 0.730 3.040 1.075 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  1.885 0.730 2.115 2.410 ;
        RECT  1.885 2.180 2.585 2.410 ;
        RECT  2.340 2.180 2.585 3.525 ;
        RECT  2.240 3.185 2.585 3.525 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.045 1.950 ;
        RECT  1.520 3.245 1.860 4.105 ;
        RECT  2.815 1.720 3.045 4.105 ;
        RECT  1.520 3.765 3.045 4.105 ;
        RECT  3.270 1.355 3.595 1.670 ;
        RECT  3.275 1.355 3.595 3.015 ;
        RECT  3.275 1.880 4.605 2.220 ;
        RECT  3.275 1.880 3.605 3.015 ;
        RECT  4.745 1.240 5.185 1.585 ;
        RECT  4.935 1.240 5.185 2.220 ;
        RECT  4.935 1.880 5.275 2.220 ;
        RECT  4.745 2.640 5.085 4.250 ;
        RECT  4.745 3.910 5.445 4.250 ;
    END
END ITLX2

MACRO ITLX16
    CLASS CORE ;
    FOREIGN ITLX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.050 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.307  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 1.880 1.560 2.165 ;
        RECT  0.750 1.640 1.135 2.165 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.040 2.070 11.395 2.410 ;
        RECT  10.835 2.070 11.215 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 9.826  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  21.490 0.700 21.925 4.150 ;
        RECT  14.040 1.840 21.925 2.440 ;
        RECT  20.050 0.700 20.390 4.150 ;
        RECT  20.040 0.700 20.390 2.440 ;
        RECT  18.610 0.700 18.955 4.150 ;
        RECT  18.600 0.700 18.955 2.440 ;
        RECT  17.170 0.700 17.510 4.150 ;
        RECT  17.165 0.700 17.510 2.440 ;
        RECT  15.730 0.700 16.070 4.150 ;
        RECT  15.725 0.700 16.070 2.440 ;
        RECT  14.290 0.700 14.640 2.440 ;
        RECT  14.290 0.700 14.630 4.150 ;
        RECT  12.845 2.850 14.630 3.080 ;
        RECT  14.040 1.150 14.630 3.080 ;
        RECT  12.690 1.150 14.640 1.380 ;
        RECT  12.845 2.850 13.185 4.150 ;
        RECT  12.690 0.880 13.030 1.380 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 22.050 0.400 ;
        RECT  20.770 -0.400 21.110 1.570 ;
        RECT  19.330 -0.400 19.670 1.570 ;
        RECT  17.890 -0.400 18.230 1.575 ;
        RECT  16.450 -0.400 16.790 1.570 ;
        RECT  15.010 -0.400 15.350 1.570 ;
        RECT  13.475 -0.400 13.815 0.920 ;
        RECT  11.965 -0.400 12.305 1.280 ;
        RECT  10.250 -0.400 10.590 0.710 ;
        RECT  8.145 -0.400 8.485 1.510 ;
        RECT  6.705 -0.400 7.045 1.115 ;
        RECT  5.265 -0.400 5.605 1.115 ;
        RECT  2.385 -0.400 2.725 1.555 ;
        RECT  0.905 -0.400 1.245 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 22.050 5.280 ;
        RECT  20.770 2.740 21.110 5.280 ;
        RECT  19.330 2.730 19.670 5.280 ;
        RECT  17.890 2.740 18.230 5.280 ;
        RECT  16.450 2.740 16.790 5.280 ;
        RECT  15.010 2.740 15.350 5.280 ;
        RECT  13.570 3.310 13.910 5.280 ;
        RECT  12.085 2.850 12.425 5.280 ;
        RECT  10.215 3.840 10.555 5.280 ;
        RECT  8.145 3.175 8.485 5.280 ;
        RECT  6.705 3.175 7.045 5.280 ;
        RECT  5.265 3.175 5.605 5.280 ;
        RECT  2.385 3.355 2.725 5.280 ;
        RECT  0.905 2.860 1.245 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.895 2.330 2.255 2.630 ;
        RECT  0.180 2.395 2.255 2.630 ;
        RECT  1.905 2.330 2.255 2.665 ;
        RECT  0.180 0.700 0.520 4.180 ;
        RECT  9.465 1.400 11.235 1.745 ;
        RECT  5.750 2.095 7.480 2.410 ;
        RECT  5.750 2.070 7.465 2.410 ;
        RECT  9.465 1.400 9.725 2.485 ;
        RECT  7.335 2.200 9.725 2.485 ;
        RECT  9.495 1.400 9.725 3.150 ;
        RECT  9.495 2.740 9.850 3.150 ;
        RECT  9.495 2.860 11.275 3.150 ;
        RECT  3.105 0.630 4.885 0.885 ;
        RECT  8.855 0.735 9.205 1.170 ;
        RECT  8.855 0.940 11.735 1.170 ;
        RECT  4.545 0.630 4.885 1.535 ;
        RECT  5.985 0.740 6.325 1.620 ;
        RECT  1.665 1.175 2.110 1.515 ;
        RECT  4.545 1.305 5.135 1.535 ;
        RECT  7.425 0.740 7.770 1.620 ;
        RECT  4.955 1.390 7.905 1.620 ;
        RECT  7.675 1.390 7.905 1.970 ;
        RECT  11.465 0.940 11.735 1.840 ;
        RECT  1.880 1.175 2.110 2.095 ;
        RECT  8.855 0.735 9.085 1.970 ;
        RECT  7.675 1.740 9.085 1.970 ;
        RECT  11.615 1.610 13.130 1.970 ;
        RECT  1.880 1.865 3.445 2.095 ;
        RECT  3.105 0.630 3.445 2.455 ;
        RECT  3.105 2.225 4.165 2.455 ;
        RECT  3.825 2.225 4.165 3.790 ;
        RECT  3.825 1.115 4.165 1.995 ;
        RECT  3.825 1.765 4.775 1.995 ;
        RECT  11.625 2.280 13.135 2.620 ;
        RECT  4.545 1.765 4.775 4.250 ;
        RECT  4.545 2.715 9.205 2.945 ;
        RECT  0.180 2.395 1.60 2.630 ;
        RECT  7.335 2.200 8.50 2.485 ;
        RECT  8.855 0.940 10.20 1.170 ;
        RECT  4.955 1.390 6.60 1.620 ;
        RECT  4.545 2.715 8.40 2.945 ;
        RECT  3.100 2.690 3.445 3.125 ;
        RECT  1.665 2.895 3.445 3.125 ;
        RECT  11.625 2.280 11.855 3.610 ;
        RECT  8.865 3.380 11.855 3.610 ;
        RECT  1.665 2.895 2.005 3.880 ;
        RECT  3.105 2.690 3.445 4.250 ;
        RECT  8.865 2.715 9.205 4.180 ;
        RECT  5.985 2.715 6.325 4.185 ;
        RECT  7.425 2.715 7.765 4.185 ;
        RECT  4.545 2.715 4.885 4.250 ;
        RECT  3.105 4.020 4.885 4.250 ;
    END
END ITLX16

MACRO ITLX12
    CLASS CORE ;
    FOREIGN ITLX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.091  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.510 2.030 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.900  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.640 2.155 9.445 2.495 ;
        RECT  8.935 2.155 9.335 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.217  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.400 0.700 16.885 4.180 ;
        RECT  10.760 1.840 16.885 2.390 ;
        RECT  16.390 0.700 16.885 2.390 ;
        RECT  14.960 0.700 15.300 4.180 ;
        RECT  14.955 0.700 15.300 2.390 ;
        RECT  13.520 0.700 13.860 4.180 ;
        RECT  13.515 0.700 13.860 2.390 ;
        RECT  12.080 0.700 12.430 2.390 ;
        RECT  12.080 0.700 12.420 4.180 ;
        RECT  10.635 2.825 10.990 4.180 ;
        RECT  10.760 0.700 10.990 4.180 ;
        RECT  10.645 2.820 10.990 4.180 ;
        RECT  10.660 0.700 10.990 1.580 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  17.115 -0.400 17.460 1.570 ;
        RECT  15.680 -0.400 16.020 1.575 ;
        RECT  14.240 -0.400 14.580 1.570 ;
        RECT  12.800 -0.400 13.140 1.570 ;
        RECT  11.355 -0.400 11.695 1.570 ;
        RECT  9.795 -0.400 10.135 0.710 ;
        RECT  8.165 -0.400 8.505 0.765 ;
        RECT  6.685 -0.400 7.025 1.110 ;
        RECT  5.245 -0.400 5.580 1.115 ;
        RECT  2.385 -0.400 2.725 1.385 ;
        RECT  0.905 -0.400 1.245 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  17.120 2.640 17.460 5.280 ;
        RECT  15.680 2.660 16.020 5.280 ;
        RECT  14.240 2.660 14.580 5.280 ;
        RECT  12.800 2.660 13.140 5.280 ;
        RECT  11.360 2.660 11.700 5.280 ;
        RECT  9.755 3.840 10.095 5.280 ;
        RECT  8.125 3.840 8.505 5.280 ;
        RECT  6.685 3.150 7.025 5.280 ;
        RECT  5.245 3.150 5.585 5.280 ;
        RECT  2.385 3.415 2.725 5.280 ;
        RECT  0.905 2.910 1.245 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.390 2.245 2.620 ;
        RECT  1.890 2.390 2.245 2.720 ;
        RECT  0.180 0.700 0.520 3.910 ;
        RECT  8.985 1.405 9.335 1.745 ;
        RECT  8.180 1.515 9.335 1.745 ;
        RECT  6.610 2.070 8.410 2.410 ;
        RECT  8.180 1.515 8.410 3.150 ;
        RECT  8.180 2.860 9.205 3.150 ;
        RECT  3.085 0.795 4.865 1.050 ;
        RECT  8.660 0.940 10.430 1.170 ;
        RECT  7.410 0.995 8.840 1.225 ;
        RECT  4.525 0.795 4.865 1.535 ;
        RECT  5.970 0.740 6.305 1.620 ;
        RECT  1.665 1.105 2.005 1.445 ;
        RECT  4.525 1.305 5.115 1.535 ;
        RECT  7.410 0.740 7.745 1.620 ;
        RECT  4.935 1.390 7.745 1.620 ;
        RECT  1.775 1.105 2.005 2.025 ;
        RECT  10.115 0.940 10.430 1.970 ;
        RECT  1.775 1.795 3.425 2.025 ;
        RECT  3.085 0.795 3.425 2.455 ;
        RECT  3.085 2.225 4.140 2.455 ;
        RECT  3.805 2.225 4.140 3.770 ;
        RECT  3.805 1.280 4.145 1.995 ;
        RECT  3.805 1.765 4.755 1.995 ;
        RECT  9.765 2.280 10.530 2.620 ;
        RECT  4.525 1.765 4.755 4.230 ;
        RECT  4.525 2.690 7.745 2.920 ;
        RECT  1.665 2.955 3.425 3.185 ;
        RECT  9.765 2.280 10.090 3.610 ;
        RECT  7.405 3.380 10.090 3.610 ;
        RECT  1.665 2.955 2.005 3.895 ;
        RECT  3.085 2.685 3.425 4.230 ;
        RECT  5.965 2.690 6.305 4.125 ;
        RECT  7.405 2.690 7.745 4.165 ;
        RECT  4.525 2.690 4.865 4.230 ;
        RECT  3.085 4.000 4.865 4.230 ;
        RECT  0.180 2.390 1.80 2.620 ;
        RECT  4.935 1.390 6.80 1.620 ;
        RECT  4.525 2.690 6.70 2.920 ;
        RECT  7.405 3.380 9.00 3.610 ;
    END
END ITLX12

MACRO ITLX1
    CLASS CORE ;
    FOREIGN ITLX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.177  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.420 1.935 2.650 3.140 ;
        RECT  2.090 1.880 2.595 2.110 ;
        RECT  2.015 2.910 2.430 4.180 ;
        RECT  2.090 1.290 2.430 2.110 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.785  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.000 1.570 3.655 2.020 ;
        RECT  3.000 1.570 3.340 2.220 ;
        RECT  2.780 0.830 3.010 1.740 ;
        RECT  2.845 1.570 3.655 1.800 ;
        RECT  1.470 0.830 3.010 1.060 ;
        RECT  1.470 0.830 1.700 2.110 ;
        RECT  1.180 1.880 1.520 2.220 ;
        END
    END A
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.691  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.450 2.190 2.680 ;
        RECT  1.850 2.340 2.190 2.680 ;
        RECT  1.435 2.450 1.765 3.240 ;
        RECT  1.410 2.450 1.765 3.215 ;
        RECT  0.575 2.450 0.915 2.790 ;
        END
    END EN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.240 2.860 3.580 5.280 ;
        RECT  0.940 3.420 1.280 5.280 ;
        RECT  0.940 3.390 1.260 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.240 -0.400 3.580 1.340 ;
        RECT  0.900 -0.400 1.240 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.700 ;
        RECT  0.115 0.630 0.345 3.380 ;
        RECT  0.115 3.035 0.520 3.380 ;
    END
END ITLX1

MACRO ITLX0
    CLASS CORE ;
    FOREIGN ITLX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.223  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.375 2.070 3.715 ;
        RECT  0.125 3.310 0.660 3.715 ;
        RECT  0.125 3.310 0.505 3.850 ;
        END
    END EN
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.471  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.970 1.740 2.310 3.135 ;
        RECT  1.280 1.740 2.310 2.020 ;
        RECT  1.280 1.510 1.765 2.020 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.148  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 0.630 2.395 1.410 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.980 3.945 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.510 -0.400 0.880 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.445 1.170 1.050 1.510 ;
        RECT  0.760 1.170 1.050 3.045 ;
        RECT  0.175 2.705 1.050 3.045 ;
    END
END ITLX0

MACRO ITLCX8
    CLASS CORE ;
    FOREIGN ITLCX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.949  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.375 1.765 11.215 2.265 ;
        RECT  10.820 0.700 11.215 2.265 ;
        RECT  10.055 1.765 10.395 3.450 ;
        RECT  9.380 0.700 9.720 2.265 ;
        RECT  8.715 1.765 9.055 3.450 ;
        RECT  7.940 0.700 8.280 2.265 ;
        RECT  7.375 1.765 7.715 3.450 ;
        RECT  7.375 1.270 7.660 3.450 ;
        RECT  6.035 2.790 7.715 3.110 ;
        RECT  6.500 1.270 7.660 1.500 ;
        RECT  6.500 0.700 6.840 1.500 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.747  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.545 4.080 2.020 ;
        RECT  1.815 1.545 4.080 1.885 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.710 0.640 2.060 ;
        RECT  0.115 1.635 0.505 2.060 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.775 2.640 11.115 5.280 ;
        RECT  9.385 3.645 9.725 5.280 ;
        RECT  8.045 3.640 8.385 5.280 ;
        RECT  6.705 3.680 7.045 5.280 ;
        RECT  4.275 3.850 4.615 5.280 ;
        RECT  2.755 4.070 3.095 5.280 ;
        RECT  0.940 3.910 1.775 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.100 -0.400 10.440 1.535 ;
        RECT  8.660 -0.400 9.000 1.535 ;
        RECT  7.220 -0.400 7.560 1.040 ;
        RECT  5.780 -0.400 6.120 1.275 ;
        RECT  4.060 -0.400 4.400 0.710 ;
        RECT  2.110 -0.400 2.450 1.315 ;
        RECT  0.650 -0.400 0.990 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.350 0.905 1.690 1.245 ;
        RECT  1.350 2.120 2.775 2.460 ;
        RECT  1.350 0.905 1.585 3.110 ;
        RECT  0.875 2.770 1.585 3.110 ;
        RECT  0.650 1.170 1.120 1.455 ;
        RECT  0.675 1.170 1.120 1.480 ;
        RECT  0.870 1.170 1.120 2.540 ;
        RECT  0.395 2.290 1.120 2.540 ;
        RECT  0.395 2.290 0.645 3.680 ;
        RECT  0.180 3.430 4.045 3.680 ;
        RECT  0.180 3.430 0.520 4.140 ;
        RECT  3.705 3.430 4.045 4.190 ;
        RECT  3.360 0.955 4.710 1.295 ;
        RECT  2.195 2.860 4.710 3.200 ;
        RECT  4.410 0.955 4.710 3.620 ;
        RECT  4.410 3.340 5.965 3.620 ;
        RECT  5.625 3.340 5.965 4.250 ;
        RECT  4.940 0.700 5.280 2.070 ;
        RECT  4.940 1.730 7.070 2.070 ;
        RECT  5.265 1.730 5.605 3.110 ;
        RECT  0.180 3.430 3.60 3.680 ;
        RECT  2.195 2.860 3.50 3.200 ;
        RECT  4.940 1.730 6.60 2.070 ;
    END
END ITLCX8

MACRO ITLCX6
    CLASS CORE ;
    FOREIGN ITLCX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.004  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.135 1.830 9.325 2.170 ;
        RECT  8.930 0.700 9.325 2.170 ;
        RECT  8.210 1.830 8.550 4.190 ;
        RECT  7.490 0.700 7.830 2.170 ;
        RECT  6.770 1.830 7.110 4.170 ;
        RECT  5.335 2.380 6.390 2.670 ;
        RECT  6.135 0.700 6.390 2.670 ;
        RECT  6.050 0.700 6.390 1.580 ;
        RECT  5.330 3.830 5.670 4.170 ;
        RECT  5.335 2.380 5.670 4.170 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.614  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.765 2.085 ;
        RECT  1.655 1.640 3.765 1.890 ;
        RECT  1.655 1.640 1.940 2.220 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.110 0.505 2.735 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.930 2.640 9.270 5.280 ;
        RECT  7.490 2.640 7.830 5.280 ;
        RECT  6.050 2.900 6.390 5.280 ;
        RECT  4.565 3.830 4.905 5.280 ;
        RECT  3.245 2.805 3.580 5.280 ;
        RECT  1.640 3.460 1.980 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.210 -0.400 8.550 1.580 ;
        RECT  6.770 -0.400 7.110 1.580 ;
        RECT  5.330 -0.400 5.670 1.510 ;
        RECT  3.550 -0.400 3.890 0.710 ;
        RECT  1.815 -0.400 2.120 0.970 ;
        RECT  0.180 -0.400 0.470 0.675 ;
        RECT  0.180 -0.400 0.465 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.695 0.725 1.585 0.990 ;
        RECT  1.245 0.630 1.585 0.990 ;
        RECT  0.295 1.170 0.890 1.510 ;
        RECT  0.635 0.865 0.890 1.910 ;
        RECT  0.625 1.170 0.890 1.910 ;
        RECT  0.735 1.730 0.965 4.140 ;
        RECT  0.735 3.800 1.125 4.140 ;
        RECT  1.120 1.220 1.460 1.515 ;
        RECT  1.120 1.220 1.445 1.545 ;
        RECT  1.120 1.220 1.425 1.550 ;
        RECT  1.195 1.220 1.425 3.020 ;
        RECT  2.270 2.120 2.555 3.020 ;
        RECT  1.195 2.680 2.555 3.020 ;
        RECT  3.050 1.070 4.230 1.410 ;
        RECT  2.785 2.315 4.230 2.575 ;
        RECT  3.995 1.070 4.230 3.600 ;
        RECT  3.990 2.315 4.230 3.600 ;
        RECT  3.990 3.260 5.105 3.600 ;
        RECT  2.785 2.315 3.015 4.180 ;
        RECT  2.515 3.320 3.015 4.180 ;
        RECT  4.460 1.810 5.905 2.150 ;
        RECT  4.460 0.700 4.800 3.030 ;
    END
END ITLCX6

MACRO ITLCX4
    CLASS CORE ;
    FOREIGN ITLCX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.642  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.770 1.970 8.065 2.305 ;
        RECT  7.670 0.700 8.065 2.305 ;
        RECT  6.950 1.970 7.290 4.180 ;
        RECT  6.230 0.700 6.570 2.305 ;
        RECT  5.510 3.740 6.000 4.080 ;
        RECT  5.770 1.970 6.000 4.080 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.330 1.710 4.320 2.050 ;
        RECT  3.330 0.630 3.560 2.050 ;
        RECT  1.365 0.630 3.560 0.860 ;
        RECT  1.365 2.250 1.765 2.630 ;
        RECT  1.365 0.630 1.595 2.630 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.660 1.930 1.135 2.270 ;
        RECT  0.750 1.600 1.135 2.270 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.670 2.640 8.010 5.280 ;
        RECT  6.230 2.640 6.570 5.280 ;
        RECT  4.790 3.740 5.130 5.280 ;
        RECT  3.430 2.810 3.775 5.280 ;
        RECT  1.990 3.370 2.330 5.280 ;
        RECT  0.900 3.800 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.950 -0.400 7.290 1.685 ;
        RECT  5.510 -0.400 5.850 1.685 ;
        RECT  3.790 -0.400 4.130 1.430 ;
        RECT  0.780 -0.400 1.120 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.630 0.520 1.700 ;
        RECT  0.165 0.630 0.430 4.140 ;
        RECT  0.165 3.800 0.520 4.140 ;
        RECT  1.825 1.360 2.265 1.700 ;
        RECT  2.035 1.360 2.265 3.140 ;
        RECT  2.035 1.980 2.375 3.140 ;
        RECT  1.125 2.860 2.375 3.140 ;
        RECT  1.125 2.860 1.465 3.200 ;
        RECT  4.630 1.110 4.970 2.670 ;
        RECT  4.630 2.330 5.485 2.670 ;
        RECT  4.630 1.110 4.920 3.000 ;
        RECT  2.495 1.090 3.050 1.430 ;
        RECT  2.710 2.280 4.400 2.580 ;
        RECT  4.100 2.280 4.400 3.490 ;
        RECT  5.150 3.000 5.490 3.490 ;
        RECT  4.100 3.230 5.490 3.490 ;
        RECT  2.710 1.090 3.050 4.180 ;
    END
END ITLCX4

MACRO ITLCX20
    CLASS CORE ;
    FOREIGN ITLCX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.279  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 0.700 20.035 3.370 ;
        RECT  10.180 1.850 20.035 2.500 ;
        RECT  18.280 1.850 18.620 3.370 ;
        RECT  18.200 0.700 18.540 2.500 ;
        RECT  17.000 1.850 17.340 3.370 ;
        RECT  16.760 0.700 17.100 2.500 ;
        RECT  15.720 1.850 16.060 3.370 ;
        RECT  15.320 0.700 15.660 2.500 ;
        RECT  14.420 1.850 14.760 3.370 ;
        RECT  13.880 0.700 14.220 2.500 ;
        RECT  13.060 1.850 13.400 4.180 ;
        RECT  12.440 0.700 12.780 2.500 ;
        RECT  11.620 1.850 11.960 4.180 ;
        RECT  11.000 0.700 11.340 2.500 ;
        RECT  10.180 1.270 10.520 4.180 ;
        RECT  8.740 2.370 10.520 2.670 ;
        RECT  8.125 1.270 10.520 1.560 ;
        RECT  9.560 0.700 9.900 1.560 ;
        RECT  8.740 2.370 9.080 4.185 ;
        RECT  8.125 0.700 8.460 1.560 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.760 2.220 ;
        END
    END A
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.276  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.640 2.450 6.810 2.700 ;
        RECT  6.425 2.240 6.810 2.700 ;
        RECT  3.640 1.805 3.980 2.700 ;
        END
    END EN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  18.920 3.590 19.260 5.280 ;
        RECT  17.640 3.595 17.980 5.280 ;
        RECT  16.360 3.595 16.700 5.280 ;
        RECT  15.070 3.580 15.410 5.280 ;
        RECT  13.780 3.590 14.120 5.280 ;
        RECT  12.340 2.730 12.680 5.280 ;
        RECT  10.900 2.730 11.240 5.280 ;
        RECT  9.460 2.900 9.800 5.280 ;
        RECT  8.070 2.690 8.360 5.280 ;
        RECT  5.860 4.080 7.270 5.280 ;
        RECT  4.380 3.390 4.720 5.280 ;
        RECT  2.940 3.390 3.280 5.280 ;
        RECT  0.900 2.960 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.620 ;
        RECT  17.480 -0.400 17.820 1.620 ;
        RECT  16.040 -0.400 16.380 1.620 ;
        RECT  14.600 -0.400 14.940 1.620 ;
        RECT  13.160 -0.400 13.500 1.620 ;
        RECT  11.720 -0.400 12.060 1.620 ;
        RECT  10.280 -0.400 10.620 1.040 ;
        RECT  8.840 -0.400 9.180 1.040 ;
        RECT  6.050 -0.400 7.510 0.655 ;
        RECT  4.180 -0.400 4.520 0.655 ;
        RECT  2.360 -0.400 2.700 0.655 ;
        RECT  0.940 -0.400 1.280 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.070 1.290 1.410 ;
        RECT  0.990 2.015 1.430 2.355 ;
        RECT  0.990 1.070 1.290 2.730 ;
        RECT  0.180 2.450 1.290 2.730 ;
        RECT  0.180 2.450 0.520 4.090 ;
        RECT  5.705 1.345 7.270 1.685 ;
        RECT  5.705 1.345 6.040 2.220 ;
        RECT  7.040 1.345 7.270 3.270 ;
        RECT  6.410 2.930 7.270 3.270 ;
        RECT  3.180 1.345 5.060 1.575 ;
        RECT  4.720 1.345 5.060 1.685 ;
        RECT  3.180 1.345 3.410 3.160 ;
        RECT  3.180 2.930 5.440 3.160 ;
        RECT  5.100 3.500 7.840 3.805 ;
        RECT  3.660 2.930 4.000 4.180 ;
        RECT  5.100 2.930 5.440 4.180 ;
        RECT  7.500 2.500 7.840 4.250 ;
        RECT  3.270 0.775 3.650 1.115 ;
        RECT  1.650 0.885 7.895 1.115 ;
        RECT  1.650 0.885 2.090 1.590 ;
        RECT  7.665 0.885 7.895 2.140 ;
        RECT  7.665 1.790 9.630 2.140 ;
        RECT  1.750 0.885 2.090 3.740 ;
        RECT  3.180 2.930 4.60 3.160 ;
        RECT  5.100 3.500 6.30 3.805 ;
        RECT  1.650 0.885 6.20 1.115 ;
    END
END ITLCX20

MACRO ITLCX16
    CLASS CORE ;
    FOREIGN ITLCX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 10.310  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 0.700 17.515 4.180 ;
        RECT  9.920 1.830 17.515 2.430 ;
        RECT  15.680 0.700 16.020 4.180 ;
        RECT  14.240 0.700 14.580 4.180 ;
        RECT  12.800 0.700 13.140 4.180 ;
        RECT  11.360 0.700 11.700 4.180 ;
        RECT  9.920 0.700 10.260 4.180 ;
        RECT  7.140 2.390 10.260 2.670 ;
        RECT  8.480 1.360 10.260 1.590 ;
        RECT  8.480 2.390 8.820 4.180 ;
        RECT  8.480 0.700 8.820 1.590 ;
        RECT  7.140 2.390 7.430 3.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.242  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.770 1.640 4.285 2.030 ;
        RECT  1.740 2.450 4.070 2.750 ;
        RECT  3.770 1.640 4.070 2.750 ;
        RECT  1.740 2.120 2.080 2.750 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.515 0.505 2.145 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.400 2.660 16.740 5.280 ;
        RECT  14.960 2.660 15.300 5.280 ;
        RECT  13.520 2.660 13.860 5.280 ;
        RECT  12.080 2.660 12.420 5.280 ;
        RECT  10.640 2.660 10.980 5.280 ;
        RECT  9.200 2.900 9.540 5.280 ;
        RECT  7.760 3.370 8.100 5.280 ;
        RECT  5.060 3.910 5.400 5.280 ;
        RECT  3.540 3.600 3.880 5.280 ;
        RECT  0.940 3.830 2.440 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.600 ;
        RECT  14.960 -0.400 15.300 1.600 ;
        RECT  13.520 -0.400 13.860 1.600 ;
        RECT  12.080 -0.400 12.420 1.600 ;
        RECT  10.640 -0.400 10.980 1.600 ;
        RECT  9.200 -0.400 9.540 1.130 ;
        RECT  7.760 -0.400 8.100 1.320 ;
        RECT  5.880 -0.400 6.220 1.305 ;
        RECT  3.960 -0.400 4.300 0.710 ;
        RECT  0.940 -0.400 2.490 0.670 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.230 1.360 2.770 1.700 ;
        RECT  2.470 1.360 2.770 2.220 ;
        RECT  1.230 1.360 1.510 3.320 ;
        RECT  1.230 2.980 1.840 3.320 ;
        RECT  0.180 0.900 3.230 1.130 ;
        RECT  0.180 0.900 1.000 1.240 ;
        RECT  3.000 0.900 3.230 2.220 ;
        RECT  3.000 1.880 3.480 2.220 ;
        RECT  0.735 0.900 1.000 2.940 ;
        RECT  0.175 2.640 1.000 2.940 ;
        RECT  0.175 2.640 0.520 3.560 ;
        RECT  3.460 1.070 4.745 1.410 ;
        RECT  2.820 3.080 4.745 3.370 ;
        RECT  4.515 1.070 4.745 3.680 ;
        RECT  4.300 2.640 4.745 3.680 ;
        RECT  4.300 3.400 6.910 3.680 ;
        RECT  2.820 3.080 3.160 4.180 ;
        RECT  6.570 2.970 6.910 4.250 ;
        RECT  4.975 0.965 5.280 2.110 ;
        RECT  6.820 0.965 7.160 2.120 ;
        RECT  4.975 1.820 9.350 2.110 ;
        RECT  6.050 1.820 9.350 2.120 ;
        RECT  6.050 1.820 6.340 3.170 ;
        RECT  0.180 0.900 2.40 1.130 ;
        RECT  4.300 3.400 5.80 3.680 ;
        RECT  4.975 1.820 8.40 2.110 ;
        RECT  6.050 1.820 8.90 2.120 ;
    END
END ITLCX16

MACRO ITLCX12
    CLASS CORE ;
    FOREIGN ITLCX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.340 1.640 13.735 4.180 ;
        RECT  7.935 1.830 13.735 2.380 ;
        RECT  12.620 1.640 13.735 2.380 ;
        RECT  12.620 0.700 12.960 2.380 ;
        RECT  11.950 1.830 12.290 3.430 ;
        RECT  11.180 0.700 11.520 2.380 ;
        RECT  10.610 1.830 10.950 3.430 ;
        RECT  9.740 0.700 10.080 2.380 ;
        RECT  9.270 1.830 9.610 3.430 ;
        RECT  7.935 1.270 8.640 2.380 ;
        RECT  8.300 0.700 8.640 2.380 ;
        RECT  7.935 1.270 8.270 3.430 ;
        RECT  6.550 2.830 8.270 3.170 ;
        RECT  6.860 1.270 8.640 1.540 ;
        RECT  6.860 0.700 7.200 1.540 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.931  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.850 2.210 4.380 2.440 ;
        RECT  3.905 1.640 4.380 2.440 ;
        RECT  1.850 2.120 2.190 2.460 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.640 0.625 2.125 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.620 3.620 12.960 5.280 ;
        RECT  11.280 3.620 11.620 5.280 ;
        RECT  9.940 3.620 10.280 5.280 ;
        RECT  8.600 3.630 8.940 5.280 ;
        RECT  7.270 3.630 7.610 5.280 ;
        RECT  4.840 3.910 5.180 5.280 ;
        RECT  3.320 4.170 3.660 5.280 ;
        RECT  2.200 4.170 2.540 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.340 -0.400 13.680 1.310 ;
        RECT  11.900 -0.400 12.240 1.580 ;
        RECT  10.460 -0.400 10.800 1.580 ;
        RECT  9.020 -0.400 9.360 1.580 ;
        RECT  7.580 -0.400 7.920 1.040 ;
        RECT  6.140 -0.400 6.480 1.540 ;
        RECT  4.360 -0.400 4.700 0.710 ;
        RECT  2.620 -0.400 2.960 1.410 ;
        RECT  0.180 -0.400 0.520 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.860 0.700 2.200 1.890 ;
        RECT  1.390 1.640 3.260 1.890 ;
        RECT  2.920 1.640 3.260 1.980 ;
        RECT  1.390 1.640 1.620 3.450 ;
        RECT  1.390 3.110 1.780 3.450 ;
        RECT  0.855 1.070 1.240 1.410 ;
        RECT  0.740 2.640 1.130 3.560 ;
        RECT  0.855 1.070 1.130 3.940 ;
        RECT  0.855 3.680 4.230 3.940 ;
        RECT  3.890 3.680 4.230 4.250 ;
        RECT  3.850 1.070 4.915 1.410 ;
        RECT  4.615 1.070 4.915 2.970 ;
        RECT  2.760 2.670 5.600 2.970 ;
        RECT  5.300 2.670 5.600 3.680 ;
        RECT  2.760 2.670 3.100 3.450 ;
        RECT  4.080 2.670 4.420 3.450 ;
        RECT  5.300 3.400 6.530 3.680 ;
        RECT  6.190 3.400 6.530 4.250 ;
        RECT  5.270 0.700 5.610 2.110 ;
        RECT  5.270 1.770 7.310 2.110 ;
        RECT  5.830 1.770 6.170 3.110 ;
        RECT  0.855 3.680 3.50 3.940 ;
        RECT  2.760 2.670 4.60 2.970 ;
        RECT  5.270 1.770 6.80 2.110 ;
    END
END ITLCX12

MACRO ITHX8
    CLASS CORE ;
    FOREIGN ITHX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.720  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.930 2.250 6.805 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 5.573  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.075 0.700 12.475 4.180 ;
        RECT  7.750 1.870 12.475 2.370 ;
        RECT  12.070 0.700 12.475 2.370 ;
        RECT  10.635 0.700 10.980 2.370 ;
        RECT  10.635 0.700 10.975 4.180 ;
        RECT  9.195 0.700 9.545 2.370 ;
        RECT  9.195 0.700 9.535 4.180 ;
        RECT  7.750 0.700 8.090 4.180 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.761  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.680 4.080 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.360 -0.400 11.700 1.600 ;
        RECT  9.920 -0.400 10.260 1.600 ;
        RECT  8.475 -0.400 8.815 1.600 ;
        RECT  6.950 -0.400 7.290 0.940 ;
        RECT  5.245 -0.400 5.585 1.020 ;
        RECT  3.805 -0.400 4.145 1.075 ;
        RECT  0.945 -0.400 1.285 1.570 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.355 2.640 11.695 5.280 ;
        RECT  9.915 2.640 10.255 5.280 ;
        RECT  8.470 2.640 8.810 5.280 ;
        RECT  6.935 3.840 7.275 5.280 ;
        RECT  5.335 3.840 5.700 5.280 ;
        RECT  3.900 3.260 4.240 5.280 ;
        RECT  0.940 2.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.800 1.435 2.140 ;
        RECT  0.180 1.175 0.520 3.220 ;
        RECT  6.105 1.635 6.445 1.970 ;
        RECT  5.345 1.740 6.445 1.970 ;
        RECT  5.345 1.740 5.580 2.410 ;
        RECT  4.320 2.070 5.580 2.410 ;
        RECT  5.350 1.740 5.580 3.150 ;
        RECT  5.350 2.865 6.450 3.150 ;
        RECT  2.385 1.150 2.725 1.995 ;
        RECT  2.385 1.765 3.410 1.995 ;
        RECT  3.180 1.765 3.410 4.250 ;
        RECT  3.180 2.640 4.980 2.870 ;
        RECT  4.620 2.640 4.980 3.610 ;
        RECT  7.190 2.310 7.520 3.610 ;
        RECT  4.620 3.380 7.520 3.610 ;
        RECT  1.660 2.685 2.000 4.250 ;
        RECT  4.620 2.640 4.960 4.185 ;
        RECT  3.180 2.640 3.520 4.250 ;
        RECT  1.660 4.020 3.520 4.250 ;
        RECT  1.665 0.630 3.425 0.885 ;
        RECT  4.525 0.700 4.865 1.650 ;
        RECT  3.085 0.630 3.425 1.535 ;
        RECT  4.525 1.250 7.520 1.405 ;
        RECT  5.760 1.170 7.520 1.405 ;
        RECT  3.085 1.305 5.930 1.480 ;
        RECT  3.085 1.305 4.870 1.535 ;
        RECT  4.525 1.250 4.870 1.650 ;
        RECT  7.225 1.170 7.520 1.980 ;
        RECT  1.665 0.630 2.005 2.455 ;
        RECT  1.665 2.225 2.720 2.455 ;
        RECT  2.380 2.225 2.720 3.790 ;
        RECT  4.620 3.380 6.50 3.610 ;
        RECT  4.525 1.250 6.70 1.405 ;
        RECT  3.085 1.305 4.70 1.480 ;
    END
END ITHX8

MACRO ITHX6
    CLASS CORE ;
    FOREIGN ITHX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.055 6.325 2.340 ;
        RECT  5.795 2.055 6.210 2.580 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.180 0.700 10.585 4.180 ;
        RECT  7.300 1.870 10.585 2.210 ;
        RECT  10.175 0.700 10.585 2.210 ;
        RECT  8.740 0.700 9.085 2.210 ;
        RECT  8.740 0.700 9.080 4.180 ;
        RECT  7.300 0.700 7.650 2.210 ;
        RECT  7.300 0.700 7.640 4.180 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.513  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.135 2.890 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.460 2.740 9.800 5.280 ;
        RECT  8.020 2.740 8.360 5.280 ;
        RECT  6.580 2.730 6.920 5.280 ;
        RECT  5.120 3.270 5.460 5.280 ;
        RECT  3.680 3.255 4.020 5.280 ;
        RECT  0.760 3.940 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.465 -0.400 9.805 1.575 ;
        RECT  8.025 -0.400 8.365 1.570 ;
        RECT  6.580 -0.400 6.920 1.365 ;
        RECT  3.825 -0.400 5.125 0.975 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.610 1.595 1.950 ;
        RECT  1.365 1.610 1.595 2.940 ;
        RECT  1.365 2.595 2.230 2.940 ;
        RECT  0.180 1.090 0.520 3.440 ;
        RECT  2.380 1.360 2.720 1.905 ;
        RECT  2.380 1.675 3.150 1.905 ;
        RECT  2.920 1.675 3.150 4.130 ;
        RECT  2.920 2.795 4.740 3.025 ;
        RECT  1.520 3.195 1.860 4.130 ;
        RECT  4.400 2.795 4.740 3.880 ;
        RECT  2.920 2.660 3.300 4.130 ;
        RECT  1.520 3.790 3.300 4.130 ;
        RECT  4.155 2.205 5.525 2.545 ;
        RECT  5.275 2.205 5.525 3.040 ;
        RECT  5.275 2.810 6.160 3.040 ;
        RECT  5.820 2.810 6.160 3.880 ;
        RECT  5.330 1.080 6.205 1.365 ;
        RECT  1.620 0.900 3.595 1.130 ;
        RECT  1.620 0.900 2.115 1.240 ;
        RECT  3.365 0.900 3.595 1.580 ;
        RECT  3.380 1.350 5.100 1.695 ;
        RECT  4.850 1.595 7.070 1.825 ;
        RECT  6.760 1.595 7.070 2.100 ;
        RECT  1.885 0.900 2.115 2.365 ;
        RECT  1.885 2.135 2.690 2.365 ;
        RECT  2.460 2.135 2.690 3.515 ;
        RECT  2.240 3.170 2.690 3.515 ;
        RECT  4.850 1.595 6.30 1.825 ;
    END
END ITHX6

MACRO ITHX4
    CLASS CORE ;
    FOREIGN ITHX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.356  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.795 2.165 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.575 0.995 8.065 4.120 ;
        RECT  6.135 1.840 8.065 2.180 ;
        RECT  6.135 0.995 6.485 2.180 ;
        RECT  6.135 0.995 6.475 4.120 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.135 2.890 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.295 2.800 8.635 5.280 ;
        RECT  6.855 2.800 7.195 5.280 ;
        RECT  5.415 2.800 5.755 5.280 ;
        RECT  3.935 2.855 5.755 3.085 ;
        RECT  3.935 2.855 4.275 3.790 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.300 -0.400 8.640 1.335 ;
        RECT  6.860 -0.400 7.200 1.335 ;
        RECT  5.415 -0.400 5.755 1.435 ;
        RECT  3.900 -0.400 4.240 0.950 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.050 2.985 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.540 0.785 2.960 1.125 ;
        RECT  1.885 0.785 2.960 1.130 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.570 2.410 ;
        RECT  2.280 2.180 2.570 3.515 ;
        RECT  3.190 1.050 3.480 1.410 ;
        RECT  3.190 1.180 4.255 1.410 ;
        RECT  4.025 1.880 4.515 2.220 ;
        RECT  4.025 1.180 4.255 2.625 ;
        RECT  3.260 2.395 4.255 2.625 ;
        RECT  3.260 2.395 3.555 3.790 ;
        RECT  2.345 1.360 2.640 1.950 ;
        RECT  2.345 1.720 3.030 1.950 ;
        RECT  1.520 3.245 1.860 4.085 ;
        RECT  2.800 1.720 3.030 4.250 ;
        RECT  1.520 3.745 3.030 4.085 ;
        RECT  4.655 3.315 4.995 4.250 ;
        RECT  2.800 4.020 4.995 4.250 ;
        RECT  4.660 1.105 5.000 1.450 ;
        RECT  4.750 1.105 5.000 2.110 ;
        RECT  4.750 1.880 5.905 2.110 ;
        RECT  5.570 1.880 5.905 2.220 ;
        RECT  2.800 4.020 3.20 4.250 ;
    END
END ITHX4

MACRO ITHX3
    CLASS CORE ;
    FOREIGN ITHX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.460 3.755 4.085 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.625 2.250 8.065 2.630 ;
        RECT  7.625 0.995 7.970 3.965 ;
        RECT  6.185 1.840 7.970 2.180 ;
        RECT  6.185 0.995 6.535 2.180 ;
        RECT  6.185 0.995 6.525 3.965 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.135 2.890 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.905 2.645 7.245 5.280 ;
        RECT  5.425 2.520 5.805 5.280 ;
        RECT  3.985 2.520 4.325 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.910 -0.400 7.250 1.335 ;
        RECT  5.465 -0.400 5.805 1.335 ;
        RECT  3.985 -0.400 4.325 1.390 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.050 2.985 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.880 0.785 3.040 1.130 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.585 2.410 ;
        RECT  2.280 2.180 2.585 3.255 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.045 1.950 ;
        RECT  1.520 3.245 1.860 3.825 ;
        RECT  2.815 1.720 3.045 3.825 ;
        RECT  1.520 3.485 3.045 3.825 ;
        RECT  3.275 1.870 4.565 2.210 ;
        RECT  3.275 1.020 3.605 3.125 ;
        RECT  4.705 2.520 5.045 4.250 ;
        RECT  4.705 1.105 5.045 1.450 ;
        RECT  4.795 1.105 5.045 2.040 ;
        RECT  4.795 1.700 5.955 2.040 ;
    END
END ITHX3

MACRO ITHX20
    CLASS CORE ;
    FOREIGN ITHX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.720 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.667  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.285 2.070 14.030 2.410 ;
        RECT  13.350 2.070 13.745 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  27.200 0.700 27.595 4.180 ;
        RECT  16.810 1.840 27.595 2.490 ;
        RECT  25.760 0.700 26.100 4.180 ;
        RECT  25.750 0.700 26.100 2.490 ;
        RECT  24.320 0.700 24.665 4.180 ;
        RECT  24.310 0.700 24.665 2.490 ;
        RECT  22.880 0.700 23.220 4.180 ;
        RECT  22.875 0.700 23.220 2.490 ;
        RECT  21.440 0.700 21.780 4.180 ;
        RECT  21.435 0.700 21.780 2.490 ;
        RECT  20.000 0.700 20.350 2.490 ;
        RECT  20.000 0.700 20.340 4.180 ;
        RECT  18.560 0.700 18.900 4.180 ;
        RECT  17.120 0.700 17.460 4.180 ;
        RECT  15.680 2.810 17.460 3.090 ;
        RECT  16.810 1.155 17.460 3.090 ;
        RECT  15.600 1.155 17.460 1.385 ;
        RECT  15.680 2.810 16.020 4.180 ;
        RECT  15.600 0.850 15.940 1.385 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.721  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.880 0.530 2.630 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 27.720 0.400 ;
        RECT  26.480 -0.400 26.820 1.570 ;
        RECT  25.040 -0.400 25.380 1.570 ;
        RECT  23.600 -0.400 23.940 1.575 ;
        RECT  22.160 -0.400 22.500 1.570 ;
        RECT  20.720 -0.400 21.060 1.570 ;
        RECT  19.280 -0.400 19.620 1.570 ;
        RECT  17.840 -0.400 18.180 1.570 ;
        RECT  16.355 -0.400 16.700 0.925 ;
        RECT  14.765 -0.400 15.105 1.195 ;
        RECT  11.585 -0.400 13.245 0.655 ;
        RECT  10.260 -0.400 10.600 1.510 ;
        RECT  8.820 -0.400 9.160 1.510 ;
        RECT  7.380 -0.400 7.720 1.140 ;
        RECT  5.940 -0.400 6.280 1.075 ;
        RECT  3.060 -0.400 3.400 1.530 ;
        RECT  1.620 -0.400 1.960 1.410 ;
        RECT  0.180 -0.400 0.520 1.650 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 27.720 5.280 ;
        RECT  26.480 2.760 26.820 5.280 ;
        RECT  25.040 2.760 25.380 5.280 ;
        RECT  23.600 2.760 23.940 5.280 ;
        RECT  22.160 2.760 22.500 5.280 ;
        RECT  20.720 2.760 21.060 5.280 ;
        RECT  19.280 2.760 19.620 5.280 ;
        RECT  17.840 2.760 18.180 5.280 ;
        RECT  16.400 3.320 16.740 5.280 ;
        RECT  14.440 3.840 15.300 5.280 ;
        RECT  14.960 2.810 15.300 5.280 ;
        RECT  12.960 3.840 13.300 5.280 ;
        RECT  11.520 3.840 11.860 5.280 ;
        RECT  10.240 3.200 10.580 5.280 ;
        RECT  8.800 3.200 9.140 5.280 ;
        RECT  7.360 3.200 7.700 5.280 ;
        RECT  5.920 3.200 6.260 5.280 ;
        RECT  3.060 3.145 3.400 5.280 ;
        RECT  1.620 2.760 1.960 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.870 2.150 2.210 ;
        RECT  0.900 0.830 1.240 3.910 ;
        RECT  11.755 1.345 14.005 1.655 ;
        RECT  5.685 2.070 7.940 2.460 ;
        RECT  5.685 2.200 12.055 2.460 ;
        RECT  11.755 1.345 12.055 3.150 ;
        RECT  11.755 2.830 12.580 3.150 ;
        RECT  11.755 2.860 14.030 3.150 ;
        RECT  4.500 1.115 4.840 1.995 ;
        RECT  4.500 1.765 5.430 1.995 ;
        RECT  14.260 2.230 16.380 2.570 ;
        RECT  5.200 1.765 5.430 4.250 ;
        RECT  2.340 2.685 4.100 2.915 ;
        RECT  5.200 2.690 11.300 2.970 ;
        RECT  10.960 2.690 11.300 3.610 ;
        RECT  14.260 2.230 14.560 3.610 ;
        RECT  10.960 3.380 14.560 3.610 ;
        RECT  3.760 2.685 4.100 4.250 ;
        RECT  6.640 2.690 6.980 4.120 ;
        RECT  8.080 2.690 8.425 4.120 ;
        RECT  9.520 2.690 9.860 4.145 ;
        RECT  2.340 2.685 2.680 4.180 ;
        RECT  5.200 2.690 5.540 4.250 ;
        RECT  3.760 3.970 5.540 4.250 ;
        RECT  3.780 0.630 5.560 0.885 ;
        RECT  10.980 0.885 14.535 1.115 ;
        RECT  5.220 0.630 5.560 1.535 ;
        RECT  6.660 0.730 7.000 1.650 ;
        RECT  2.340 1.190 2.680 1.530 ;
        RECT  5.220 1.305 7.000 1.535 ;
        RECT  14.260 0.885 14.535 1.900 ;
        RECT  8.100 0.740 8.440 1.650 ;
        RECT  6.660 1.370 8.440 1.650 ;
        RECT  8.170 0.740 8.440 1.970 ;
        RECT  9.540 0.740 9.880 1.970 ;
        RECT  14.260 1.615 16.385 1.900 ;
        RECT  10.980 0.885 11.320 1.970 ;
        RECT  8.170 1.740 11.320 1.970 ;
        RECT  2.380 1.190 2.680 2.455 ;
        RECT  3.780 0.630 4.120 2.455 ;
        RECT  2.380 2.225 4.820 2.455 ;
        RECT  4.480 2.225 4.820 3.740 ;
        RECT  11.755 1.345 13.60 1.655 ;
        RECT  5.685 2.070 6.80 2.460 ;
        RECT  5.685 2.200 11.90 2.460 ;
        RECT  11.755 2.860 13.50 3.150 ;
        RECT  14.260 2.230 15.60 2.570 ;
        RECT  5.200 2.690 10.70 2.970 ;
        RECT  10.960 3.380 13.60 3.610 ;
        RECT  10.980 0.885 13.90 1.115 ;
        RECT  14.260 1.615 15.70 1.900 ;
        RECT  8.170 1.740 10.60 1.970 ;
        RECT  2.380 2.225 3.70 2.455 ;
    END
END ITHX20

MACRO ITHX2
    CLASS CORE ;
    FOREIGN ITHX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 3.460 3.760 4.085 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.084  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.945 0.995 7.435 3.965 ;
        RECT  5.505 1.840 7.435 2.180 ;
        RECT  5.505 0.995 5.855 2.180 ;
        RECT  5.505 0.995 5.845 3.680 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.135 2.890 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.225 2.645 6.565 5.280 ;
        RECT  4.025 2.640 4.365 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.230 -0.400 6.570 1.335 ;
        RECT  4.025 -0.400 4.365 1.585 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.050 2.985 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.880 0.730 3.040 1.075 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  1.885 0.730 2.115 2.410 ;
        RECT  1.885 2.180 2.585 2.410 ;
        RECT  2.280 2.180 2.585 3.255 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.045 1.950 ;
        RECT  1.520 3.245 1.860 3.825 ;
        RECT  2.815 1.720 3.045 3.825 ;
        RECT  1.520 3.485 3.045 3.825 ;
        RECT  3.270 1.355 3.595 1.670 ;
        RECT  3.275 1.355 3.595 3.015 ;
        RECT  3.275 1.880 4.605 2.220 ;
        RECT  3.275 1.880 3.605 3.015 ;
        RECT  4.745 1.240 5.275 1.585 ;
        RECT  4.835 1.240 5.275 2.220 ;
        RECT  4.745 2.640 5.085 4.250 ;
        RECT  4.745 3.910 5.445 4.250 ;
    END
END ITHX2

MACRO ITHX16
    CLASS CORE ;
    FOREIGN ITHX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.050 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.040 2.070 11.395 2.410 ;
        RECT  10.835 2.070 11.215 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 9.826  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  21.490 0.700 21.925 4.150 ;
        RECT  14.040 1.840 21.925 2.440 ;
        RECT  20.050 0.700 20.390 4.150 ;
        RECT  20.040 0.700 20.390 2.440 ;
        RECT  18.610 0.700 18.955 4.150 ;
        RECT  18.600 0.700 18.955 2.440 ;
        RECT  17.170 0.700 17.510 4.150 ;
        RECT  17.165 0.700 17.510 2.440 ;
        RECT  15.730 0.700 16.070 4.150 ;
        RECT  15.725 0.700 16.070 2.440 ;
        RECT  14.290 0.700 14.640 2.440 ;
        RECT  14.290 0.700 14.630 4.150 ;
        RECT  12.845 2.850 14.630 3.080 ;
        RECT  14.040 1.150 14.630 3.080 ;
        RECT  12.690 1.150 14.640 1.380 ;
        RECT  12.845 2.850 13.185 4.150 ;
        RECT  12.690 0.880 13.030 1.380 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.255  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 3.470 1.790 4.250 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 22.050 0.400 ;
        RECT  20.770 -0.400 21.110 1.570 ;
        RECT  19.330 -0.400 19.670 1.570 ;
        RECT  17.890 -0.400 18.230 1.575 ;
        RECT  16.450 -0.400 16.790 1.570 ;
        RECT  15.010 -0.400 15.350 1.570 ;
        RECT  13.475 -0.400 13.815 0.920 ;
        RECT  11.965 -0.400 12.305 1.280 ;
        RECT  10.260 -0.400 10.600 0.710 ;
        RECT  8.145 -0.400 8.485 1.510 ;
        RECT  6.705 -0.400 7.045 1.115 ;
        RECT  5.265 -0.400 5.605 1.115 ;
        RECT  2.385 -0.400 2.725 1.555 ;
        RECT  0.905 -0.400 1.245 1.650 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 22.050 5.280 ;
        RECT  20.770 2.740 21.110 5.280 ;
        RECT  19.330 2.730 19.670 5.280 ;
        RECT  17.890 2.740 18.230 5.280 ;
        RECT  16.450 2.740 16.790 5.280 ;
        RECT  15.010 2.740 15.350 5.280 ;
        RECT  13.570 3.310 13.910 5.280 ;
        RECT  12.085 2.850 12.425 5.280 ;
        RECT  10.215 3.840 10.555 5.280 ;
        RECT  8.145 3.175 8.485 5.280 ;
        RECT  6.705 3.175 7.045 5.280 ;
        RECT  5.265 3.175 5.605 5.280 ;
        RECT  2.385 3.145 2.725 5.280 ;
        RECT  0.905 2.690 1.245 3.030 ;
        RECT  0.905 2.690 1.205 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.880 1.435 2.220 ;
        RECT  0.180 0.700 0.520 4.180 ;
        RECT  9.465 1.400 11.235 1.745 ;
        RECT  5.750 2.095 7.480 2.410 ;
        RECT  5.750 2.070 7.465 2.410 ;
        RECT  9.465 1.400 9.810 2.485 ;
        RECT  7.335 2.200 9.810 2.485 ;
        RECT  9.495 1.400 9.810 3.150 ;
        RECT  9.495 2.740 9.850 3.150 ;
        RECT  9.495 2.860 11.275 3.150 ;
        RECT  3.105 0.630 4.885 0.885 ;
        RECT  8.855 0.735 9.205 1.170 ;
        RECT  8.855 0.940 11.735 1.170 ;
        RECT  4.545 0.630 4.885 1.535 ;
        RECT  5.985 0.740 6.325 1.620 ;
        RECT  4.545 1.305 5.135 1.535 ;
        RECT  7.425 0.740 7.770 1.620 ;
        RECT  4.955 1.390 7.905 1.620 ;
        RECT  7.675 1.390 7.905 1.970 ;
        RECT  11.465 0.940 11.735 1.840 ;
        RECT  8.855 0.735 9.085 1.970 ;
        RECT  7.675 1.740 9.085 1.970 ;
        RECT  11.615 1.610 13.130 1.970 ;
        RECT  1.665 1.215 2.005 2.455 ;
        RECT  3.105 0.630 3.445 2.455 ;
        RECT  1.665 2.225 4.165 2.455 ;
        RECT  3.825 2.225 4.165 3.790 ;
        RECT  3.825 1.115 4.165 1.995 ;
        RECT  3.825 1.765 4.775 1.995 ;
        RECT  11.625 2.280 13.135 2.620 ;
        RECT  4.545 1.765 4.775 4.250 ;
        RECT  1.665 2.685 3.445 2.915 ;
        RECT  4.545 2.715 9.205 2.945 ;
        RECT  1.665 2.685 2.005 3.240 ;
        RECT  11.625 2.280 11.855 3.610 ;
        RECT  8.865 3.380 11.855 3.610 ;
        RECT  3.105 2.685 3.445 4.250 ;
        RECT  8.865 2.715 9.205 4.180 ;
        RECT  5.985 2.715 6.325 4.185 ;
        RECT  7.425 2.715 7.765 4.185 ;
        RECT  4.545 2.715 4.885 4.250 ;
        RECT  3.105 4.020 4.885 4.250 ;
        RECT  7.335 2.200 8.60 2.485 ;
        RECT  8.855 0.940 10.80 1.170 ;
        RECT  4.955 1.390 6.30 1.620 ;
        RECT  1.665 2.225 3.40 2.455 ;
        RECT  4.545 2.715 8.60 2.945 ;
        RECT  8.865 3.380 10.70 3.610 ;
    END
END ITHX16

MACRO ITHX12
    CLASS CORE ;
    FOREIGN ITHX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.900  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.640 2.155 9.445 2.495 ;
        RECT  8.935 2.155 9.335 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.217  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.400 0.700 16.885 4.180 ;
        RECT  10.760 1.840 16.885 2.390 ;
        RECT  16.390 0.700 16.885 2.390 ;
        RECT  14.960 0.700 15.300 4.180 ;
        RECT  14.955 0.700 15.300 2.390 ;
        RECT  13.520 0.700 13.860 4.180 ;
        RECT  13.515 0.700 13.860 2.390 ;
        RECT  12.080 0.700 12.430 2.390 ;
        RECT  12.080 0.700 12.420 4.180 ;
        RECT  10.635 2.825 10.990 4.180 ;
        RECT  10.760 0.700 10.990 4.180 ;
        RECT  10.660 0.700 10.990 1.580 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.060  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 3.470 1.790 4.250 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  17.115 -0.400 17.460 1.570 ;
        RECT  15.680 -0.400 16.020 1.575 ;
        RECT  14.240 -0.400 14.580 1.570 ;
        RECT  12.800 -0.400 13.140 1.570 ;
        RECT  11.355 -0.400 11.695 1.570 ;
        RECT  9.795 -0.400 10.135 0.710 ;
        RECT  8.165 -0.400 8.505 0.765 ;
        RECT  6.685 -0.400 7.025 1.115 ;
        RECT  5.245 -0.400 5.585 1.115 ;
        RECT  2.385 -0.400 2.725 1.570 ;
        RECT  0.905 -0.400 1.245 1.620 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  17.120 2.640 17.460 5.280 ;
        RECT  15.680 2.660 16.020 5.280 ;
        RECT  14.240 2.660 14.580 5.280 ;
        RECT  12.800 2.660 13.140 5.280 ;
        RECT  11.360 2.660 11.700 5.280 ;
        RECT  9.755 3.840 10.095 5.280 ;
        RECT  8.125 3.840 8.505 5.280 ;
        RECT  6.685 3.200 7.025 5.280 ;
        RECT  5.245 3.200 5.585 5.280 ;
        RECT  2.385 3.145 2.725 5.280 ;
        RECT  0.905 2.690 1.245 3.030 ;
        RECT  0.905 2.690 1.205 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.880 1.435 2.220 ;
        RECT  0.180 0.810 0.520 3.910 ;
        RECT  8.985 1.405 9.335 1.745 ;
        RECT  8.180 1.455 9.335 1.745 ;
        RECT  6.605 2.070 8.410 2.410 ;
        RECT  8.180 1.455 8.410 3.150 ;
        RECT  8.180 2.860 9.205 3.150 ;
        RECT  3.085 0.795 4.865 1.050 ;
        RECT  8.660 0.940 10.430 1.170 ;
        RECT  7.405 0.995 8.840 1.225 ;
        RECT  4.525 0.795 4.865 1.535 ;
        RECT  5.965 0.740 6.305 1.620 ;
        RECT  4.525 1.305 5.115 1.535 ;
        RECT  7.405 0.740 7.745 1.620 ;
        RECT  4.935 1.390 7.745 1.620 ;
        RECT  10.115 0.940 10.430 1.970 ;
        RECT  1.665 1.215 2.005 2.455 ;
        RECT  3.085 0.795 3.425 2.455 ;
        RECT  1.665 2.225 4.145 2.455 ;
        RECT  3.805 2.225 4.145 3.770 ;
        RECT  3.805 1.280 4.145 1.995 ;
        RECT  3.805 1.765 4.755 1.995 ;
        RECT  9.765 2.280 10.530 2.620 ;
        RECT  4.525 1.765 4.755 4.230 ;
        RECT  1.665 2.685 3.425 2.915 ;
        RECT  4.525 2.690 7.745 2.970 ;
        RECT  1.665 2.685 2.005 3.205 ;
        RECT  9.765 2.280 10.090 3.610 ;
        RECT  7.405 3.380 10.090 3.610 ;
        RECT  3.085 2.685 3.425 4.230 ;
        RECT  5.965 2.690 6.305 4.125 ;
        RECT  7.405 2.690 7.745 4.165 ;
        RECT  4.525 2.690 4.865 4.230 ;
        RECT  3.085 4.000 4.865 4.230 ;
        RECT  4.935 1.390 6.60 1.620 ;
        RECT  1.665 2.225 3.60 2.455 ;
        RECT  4.525 2.690 6.90 2.970 ;
        RECT  7.405 3.380 9.70 3.610 ;
    END
END ITHX12

MACRO ITHX1
    CLASS CORE ;
    FOREIGN ITHX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.177  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.420 1.935 2.650 3.140 ;
        RECT  2.090 1.880 2.595 2.110 ;
        RECT  2.015 2.910 2.430 4.180 ;
        RECT  2.090 1.290 2.430 2.110 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.785  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.000 1.570 3.655 2.020 ;
        RECT  3.000 1.570 3.340 2.220 ;
        RECT  2.780 0.830 3.010 1.740 ;
        RECT  2.845 1.570 3.655 1.800 ;
        RECT  1.515 0.830 3.010 1.060 ;
        RECT  1.515 0.830 1.745 2.110 ;
        RECT  1.180 1.880 1.520 2.220 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.469  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.660 3.950 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.240 2.860 3.580 5.280 ;
        RECT  0.940 2.910 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.240 -0.400 3.580 1.340 ;
        RECT  0.940 -0.400 1.285 1.490 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.850 2.340 2.190 2.680 ;
        RECT  0.180 2.450 2.190 2.680 ;
        RECT  0.180 1.360 0.520 3.240 ;
        RECT  0.180 2.450 1.00 2.680 ;
    END
END ITHX1

MACRO ITHX0
    CLASS CORE ;
    FOREIGN ITHX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.180  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.325 0.660 3.850 ;
        END
    END E
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.499  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 1.410 2.395 2.020 ;
        RECT  2.010 1.410 2.390 3.185 ;
        RECT  1.280 1.410 2.395 1.725 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.955 1.400 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.980 3.675 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.285 -0.400 1.095 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.175 1.170 0.785 1.510 ;
        RECT  0.175 1.170 0.405 3.095 ;
        RECT  0.175 2.755 0.520 3.095 ;
        RECT  0.175 2.860 1.780 3.095 ;
        RECT  1.550 2.860 1.780 3.765 ;
        RECT  1.550 3.425 2.070 3.765 ;
    END
END ITHX0

MACRO ITHCX8
    CLASS CORE ;
    FOREIGN ITHCX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.949  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.375 1.765 11.215 2.265 ;
        RECT  10.820 0.700 11.215 2.265 ;
        RECT  10.050 1.765 10.390 3.450 ;
        RECT  9.380 0.700 9.720 2.265 ;
        RECT  8.715 1.765 9.055 3.450 ;
        RECT  7.940 0.700 8.280 2.265 ;
        RECT  7.375 1.765 7.715 3.450 ;
        RECT  7.375 1.270 7.660 3.450 ;
        RECT  6.035 2.770 7.715 3.110 ;
        RECT  6.500 1.270 7.660 1.500 ;
        RECT  6.500 0.700 6.840 1.500 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.785  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.935 2.115 2.415 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.710 0.640 2.060 ;
        RECT  0.115 1.635 0.505 2.060 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.775 2.640 11.115 5.280 ;
        RECT  9.385 3.645 9.725 5.280 ;
        RECT  8.045 3.640 8.385 5.280 ;
        RECT  6.705 3.680 7.045 5.280 ;
        RECT  4.275 3.850 4.615 5.280 ;
        RECT  2.755 3.960 3.095 5.280 ;
        RECT  0.940 3.910 1.775 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.100 -0.400 10.440 1.535 ;
        RECT  8.660 -0.400 9.000 1.535 ;
        RECT  7.220 -0.400 7.560 1.040 ;
        RECT  5.780 -0.400 6.120 1.275 ;
        RECT  4.060 -0.400 4.400 0.710 ;
        RECT  2.110 -0.400 2.450 1.315 ;
        RECT  0.650 -0.400 0.990 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.650 1.170 1.120 1.455 ;
        RECT  0.675 1.170 1.120 1.480 ;
        RECT  0.870 1.170 1.120 2.540 ;
        RECT  0.395 2.290 1.120 2.540 ;
        RECT  0.395 2.290 0.645 3.680 ;
        RECT  0.180 3.430 4.045 3.680 ;
        RECT  3.705 3.430 4.045 4.080 ;
        RECT  0.180 3.430 0.520 4.140 ;
        RECT  1.350 1.545 4.080 1.885 ;
        RECT  1.350 0.905 1.690 3.110 ;
        RECT  0.875 2.770 1.690 3.110 ;
        RECT  3.360 0.955 4.710 1.295 ;
        RECT  2.195 2.860 4.710 3.200 ;
        RECT  4.410 0.955 4.710 3.620 ;
        RECT  4.410 3.340 5.965 3.620 ;
        RECT  5.625 3.340 5.965 4.250 ;
        RECT  4.940 0.700 5.280 2.070 ;
        RECT  4.940 1.730 7.070 2.070 ;
        RECT  5.265 1.730 5.605 3.110 ;
        RECT  0.180 3.430 3.30 3.680 ;
        RECT  1.350 1.545 3.20 1.885 ;
        RECT  2.195 2.860 3.70 3.200 ;
        RECT  4.940 1.730 6.70 2.070 ;
    END
END ITHCX8

MACRO ITHCX6
    CLASS CORE ;
    FOREIGN ITHCX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.035  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.770 1.830 9.325 2.170 ;
        RECT  8.930 0.700 9.325 2.170 ;
        RECT  8.210 1.830 8.550 4.190 ;
        RECT  7.490 0.700 7.830 2.170 ;
        RECT  6.770 1.310 7.110 4.170 ;
        RECT  5.330 2.380 7.110 2.670 ;
        RECT  6.050 1.310 7.110 1.580 ;
        RECT  6.050 0.700 6.390 1.580 ;
        RECT  5.330 2.380 5.670 4.170 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.562  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.880 1.785 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.575 2.120 1.155 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.930 2.640 9.270 5.280 ;
        RECT  7.490 2.640 7.830 5.280 ;
        RECT  6.050 2.900 6.390 5.280 ;
        RECT  4.495 3.830 4.835 5.280 ;
        RECT  3.005 2.805 3.350 5.280 ;
        RECT  1.420 3.460 1.760 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.210 -0.400 8.550 1.580 ;
        RECT  6.770 -0.400 7.110 1.080 ;
        RECT  5.330 -0.400 5.670 1.510 ;
        RECT  3.550 -0.400 3.890 0.710 ;
        RECT  1.815 -0.400 2.120 0.970 ;
        RECT  0.180 -0.400 0.490 0.685 ;
        RECT  0.180 -0.400 0.465 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.695 0.825 1.585 1.080 ;
        RECT  1.245 0.630 1.585 1.080 ;
        RECT  0.635 0.865 0.890 1.510 ;
        RECT  0.115 1.170 0.890 1.510 ;
        RECT  0.115 1.170 0.345 4.140 ;
        RECT  0.115 3.800 0.905 4.140 ;
        RECT  1.120 1.310 2.285 1.650 ;
        RECT  2.015 1.745 3.580 2.085 ;
        RECT  2.015 1.310 2.285 3.090 ;
        RECT  0.770 2.860 2.285 3.090 ;
        RECT  0.770 2.860 1.110 3.200 ;
        RECT  3.050 1.160 4.070 1.500 ;
        RECT  2.515 2.315 4.070 2.575 ;
        RECT  3.810 1.160 4.070 3.600 ;
        RECT  3.810 3.260 5.075 3.600 ;
        RECT  2.515 2.315 2.775 4.180 ;
        RECT  2.285 3.320 2.775 4.180 ;
        RECT  4.460 0.700 4.800 2.150 ;
        RECT  4.300 1.810 6.150 2.150 ;
        RECT  4.300 1.810 4.640 3.030 ;
    END
END ITHCX6

MACRO ITHCX4
    CLASS CORE ;
    FOREIGN ITHCX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.646  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.140 1.970 7.435 2.310 ;
        RECT  7.040 0.700 7.435 2.310 ;
        RECT  6.320 1.970 6.660 4.180 ;
        RECT  5.600 0.700 5.940 2.310 ;
        RECT  4.880 3.740 5.370 4.080 ;
        RECT  5.140 1.970 5.370 4.080 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.551  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 2.115 1.765 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.620 1.930 1.135 2.270 ;
        RECT  0.750 1.600 1.135 2.270 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 2.640 7.380 5.280 ;
        RECT  5.600 3.840 5.940 5.280 ;
        RECT  4.160 3.740 4.500 5.280 ;
        RECT  2.850 3.720 3.195 5.280 ;
        RECT  1.370 3.460 1.710 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.685 ;
        RECT  4.840 -0.400 5.180 0.710 ;
        RECT  3.375 -0.400 3.660 1.410 ;
        RECT  0.735 -0.400 1.080 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.505 1.700 ;
        RECT  0.115 1.335 0.520 1.700 ;
        RECT  0.115 0.630 0.390 4.180 ;
        RECT  0.115 3.840 0.735 4.180 ;
        RECT  1.470 0.630 3.145 0.860 ;
        RECT  1.470 0.630 1.810 1.885 ;
        RECT  2.915 0.630 3.145 2.050 ;
        RECT  1.470 1.655 2.225 1.885 ;
        RECT  2.915 1.710 3.850 2.050 ;
        RECT  0.810 2.715 1.150 3.090 ;
        RECT  1.995 1.655 2.225 3.090 ;
        RECT  0.810 2.860 2.225 3.090 ;
        RECT  4.160 1.190 4.500 2.690 ;
        RECT  4.160 2.350 4.905 2.690 ;
        RECT  4.040 2.370 4.345 2.970 ;
        RECT  4.040 2.370 4.340 3.000 ;
        RECT  2.080 1.140 2.685 1.425 ;
        RECT  2.455 1.140 2.685 3.490 ;
        RECT  2.455 3.230 4.910 3.490 ;
        RECT  4.570 3.020 4.910 3.490 ;
        RECT  2.130 3.320 2.620 4.180 ;
        RECT  2.455 3.230 3.60 3.490 ;
    END
END ITHCX4

MACRO ITHCX20
    CLASS CORE ;
    FOREIGN ITHCX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.279  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 0.700 20.035 3.370 ;
        RECT  10.180 1.850 20.035 2.500 ;
        RECT  18.280 1.850 18.620 3.370 ;
        RECT  18.200 0.700 18.540 2.500 ;
        RECT  17.000 1.850 17.340 3.370 ;
        RECT  16.760 0.700 17.100 2.500 ;
        RECT  15.720 1.850 16.060 3.370 ;
        RECT  15.320 0.700 15.660 2.500 ;
        RECT  14.420 1.850 14.760 3.370 ;
        RECT  13.880 0.700 14.220 2.500 ;
        RECT  13.060 1.850 13.400 4.180 ;
        RECT  12.440 0.700 12.780 2.500 ;
        RECT  11.620 1.850 11.960 4.180 ;
        RECT  11.000 0.700 11.340 2.500 ;
        RECT  10.180 1.270 10.520 4.180 ;
        RECT  8.740 2.370 10.520 2.670 ;
        RECT  8.125 1.270 10.520 1.560 ;
        RECT  9.560 0.700 9.900 1.560 ;
        RECT  8.740 2.370 9.080 4.185 ;
        RECT  8.125 0.700 8.460 1.560 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.760 2.220 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.451  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.080 6.950 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  18.920 3.610 19.260 5.280 ;
        RECT  17.640 3.615 17.980 5.280 ;
        RECT  16.360 3.615 16.700 5.280 ;
        RECT  15.070 3.615 15.410 5.280 ;
        RECT  13.780 3.625 14.120 5.280 ;
        RECT  12.340 2.730 12.680 5.280 ;
        RECT  10.900 2.730 11.240 5.280 ;
        RECT  9.460 2.900 9.800 5.280 ;
        RECT  8.070 2.690 8.360 5.280 ;
        RECT  5.860 4.170 7.270 5.280 ;
        RECT  4.380 3.165 4.720 5.280 ;
        RECT  2.940 3.165 3.280 5.280 ;
        RECT  0.900 2.960 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.620 ;
        RECT  17.480 -0.400 17.820 1.620 ;
        RECT  16.040 -0.400 16.380 1.620 ;
        RECT  14.600 -0.400 14.940 1.620 ;
        RECT  13.160 -0.400 13.500 1.620 ;
        RECT  11.720 -0.400 12.060 1.620 ;
        RECT  10.280 -0.400 10.620 1.040 ;
        RECT  8.840 -0.400 9.180 1.040 ;
        RECT  6.090 -0.400 7.550 0.655 ;
        RECT  4.220 -0.400 4.560 0.655 ;
        RECT  2.360 -0.400 2.700 0.655 ;
        RECT  0.940 -0.400 1.280 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.070 1.290 1.410 ;
        RECT  0.990 2.015 1.430 2.355 ;
        RECT  0.990 1.070 1.290 2.730 ;
        RECT  0.180 2.450 1.290 2.730 ;
        RECT  0.180 2.450 0.520 4.090 ;
        RECT  5.915 1.360 6.990 1.700 ;
        RECT  3.640 1.805 3.980 2.170 ;
        RECT  3.640 1.870 6.195 2.170 ;
        RECT  5.915 1.360 6.195 3.235 ;
        RECT  5.915 2.895 6.760 3.235 ;
        RECT  3.180 1.345 5.100 1.575 ;
        RECT  4.760 1.345 5.100 1.640 ;
        RECT  3.180 1.345 3.410 2.935 ;
        RECT  3.180 2.640 5.440 2.935 ;
        RECT  5.100 3.465 7.840 3.805 ;
        RECT  3.660 2.640 4.000 4.180 ;
        RECT  5.100 2.640 5.440 4.180 ;
        RECT  7.500 2.500 7.840 4.250 ;
        RECT  3.310 0.775 3.650 1.115 ;
        RECT  1.650 0.885 7.895 1.115 ;
        RECT  1.650 0.885 2.090 1.590 ;
        RECT  7.665 0.885 7.895 2.140 ;
        RECT  7.665 1.790 9.630 2.140 ;
        RECT  1.750 0.885 2.090 3.740 ;
        RECT  3.640 1.870 5.50 2.170 ;
        RECT  3.180 2.640 4.80 2.935 ;
        RECT  5.100 3.465 6.20 3.805 ;
        RECT  1.650 0.885 6.30 1.115 ;
    END
END ITHCX20

MACRO ITHCX16
    CLASS CORE ;
    FOREIGN ITHCX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 10.310  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 0.700 17.515 4.180 ;
        RECT  9.920 1.830 17.515 2.430 ;
        RECT  15.680 0.700 16.020 4.180 ;
        RECT  14.240 0.700 14.580 4.180 ;
        RECT  12.800 0.700 13.140 4.180 ;
        RECT  11.360 0.700 11.700 4.180 ;
        RECT  9.920 0.700 10.260 4.180 ;
        RECT  7.140 2.390 10.260 2.670 ;
        RECT  8.480 1.360 10.260 1.590 ;
        RECT  8.480 2.390 8.820 4.180 ;
        RECT  8.480 0.700 8.820 1.590 ;
        RECT  7.140 2.390 7.430 3.180 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.188  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.975 2.665 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.620 0.720 2.040 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.400 2.660 16.740 5.280 ;
        RECT  14.960 2.660 15.300 5.280 ;
        RECT  13.520 2.660 13.860 5.280 ;
        RECT  12.080 2.660 12.420 5.280 ;
        RECT  10.640 2.660 10.980 5.280 ;
        RECT  9.200 2.900 9.540 5.280 ;
        RECT  7.760 3.370 8.100 5.280 ;
        RECT  5.060 3.910 5.400 5.280 ;
        RECT  3.540 3.840 3.880 5.280 ;
        RECT  0.940 3.830 2.440 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.600 ;
        RECT  14.960 -0.400 15.300 1.600 ;
        RECT  13.520 -0.400 13.860 1.600 ;
        RECT  12.080 -0.400 12.420 1.600 ;
        RECT  10.640 -0.400 10.980 1.600 ;
        RECT  9.200 -0.400 9.540 1.130 ;
        RECT  7.760 -0.400 8.100 1.320 ;
        RECT  5.880 -0.400 6.220 1.305 ;
        RECT  3.960 -0.400 4.300 0.710 ;
        RECT  0.940 -0.400 2.490 0.670 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.900 3.125 1.130 ;
        RECT  0.180 0.900 1.230 1.240 ;
        RECT  2.895 0.900 3.125 2.460 ;
        RECT  2.895 2.120 3.480 2.460 ;
        RECT  0.950 0.900 1.230 2.940 ;
        RECT  0.175 2.640 1.230 2.940 ;
        RECT  0.175 2.640 0.520 3.560 ;
        RECT  1.500 1.360 1.840 1.700 ;
        RECT  3.840 1.690 4.280 2.030 ;
        RECT  1.500 1.360 1.785 3.195 ;
        RECT  3.840 1.690 4.070 3.090 ;
        RECT  1.500 2.860 4.070 3.090 ;
        RECT  1.500 2.860 1.840 3.195 ;
        RECT  3.420 1.120 4.740 1.460 ;
        RECT  4.300 2.640 4.740 3.610 ;
        RECT  4.510 1.120 4.740 3.610 ;
        RECT  2.820 3.320 4.740 3.610 ;
        RECT  2.820 3.330 6.910 3.610 ;
        RECT  2.820 3.320 3.160 4.180 ;
        RECT  6.570 2.970 6.910 4.250 ;
        RECT  4.970 0.965 5.280 2.110 ;
        RECT  6.820 0.965 7.160 2.120 ;
        RECT  4.970 1.820 9.350 2.110 ;
        RECT  6.050 1.820 9.350 2.120 ;
        RECT  6.050 1.820 6.340 3.100 ;
        RECT  0.180 0.900 2.20 1.130 ;
        RECT  1.500 2.860 3.50 3.090 ;
        RECT  2.820 3.330 5.10 3.610 ;
        RECT  4.970 1.820 8.40 2.110 ;
        RECT  6.050 1.820 8.80 2.120 ;
    END
END ITHCX16

MACRO ITHCX12
    CLASS CORE ;
    FOREIGN ITHCX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.340 1.640 13.735 4.180 ;
        RECT  7.935 1.830 13.735 2.380 ;
        RECT  12.620 1.640 13.735 2.380 ;
        RECT  12.620 0.700 12.960 2.380 ;
        RECT  11.950 1.830 12.290 3.430 ;
        RECT  11.180 0.700 11.520 2.380 ;
        RECT  10.610 1.830 10.950 3.430 ;
        RECT  9.740 0.700 10.080 2.380 ;
        RECT  9.270 1.830 9.610 3.430 ;
        RECT  7.935 1.270 8.640 2.380 ;
        RECT  8.300 0.700 8.640 2.380 ;
        RECT  7.935 1.270 8.270 3.430 ;
        RECT  6.550 2.830 8.270 3.170 ;
        RECT  6.860 1.270 8.640 1.540 ;
        RECT  6.860 0.700 7.200 1.540 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.955  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.635 1.860 2.150 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.640 0.625 2.125 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.620 3.620 12.960 5.280 ;
        RECT  11.280 3.620 11.620 5.280 ;
        RECT  9.940 3.620 10.280 5.280 ;
        RECT  8.600 3.630 8.940 5.280 ;
        RECT  7.270 3.630 7.610 5.280 ;
        RECT  4.840 3.910 5.180 5.280 ;
        RECT  3.320 4.170 3.660 5.280 ;
        RECT  2.200 4.170 2.540 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.340 -0.400 13.680 1.310 ;
        RECT  11.900 -0.400 12.240 1.580 ;
        RECT  10.460 -0.400 10.800 1.580 ;
        RECT  9.020 -0.400 9.360 1.580 ;
        RECT  7.580 -0.400 7.920 1.040 ;
        RECT  6.140 -0.400 6.480 1.540 ;
        RECT  4.360 -0.400 4.700 0.710 ;
        RECT  2.620 -0.400 2.960 1.460 ;
        RECT  0.180 -0.400 0.520 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.855 1.070 1.240 1.410 ;
        RECT  0.740 2.640 1.155 2.980 ;
        RECT  0.855 1.070 1.155 3.940 ;
        RECT  0.855 3.680 4.230 3.940 ;
        RECT  3.890 3.680 4.230 4.250 ;
        RECT  1.860 0.905 2.390 1.245 ;
        RECT  2.090 1.690 4.380 2.030 ;
        RECT  2.090 0.905 2.390 2.895 ;
        RECT  1.440 2.640 2.390 2.895 ;
        RECT  1.440 2.640 1.780 3.450 ;
        RECT  3.850 1.075 4.915 1.415 ;
        RECT  4.615 1.075 4.915 2.935 ;
        RECT  2.760 2.640 5.600 2.935 ;
        RECT  5.300 2.640 5.600 3.680 ;
        RECT  2.760 2.640 3.100 3.450 ;
        RECT  4.080 2.640 4.420 3.450 ;
        RECT  5.300 3.400 6.530 3.680 ;
        RECT  6.190 3.400 6.530 4.250 ;
        RECT  5.270 0.700 5.610 2.110 ;
        RECT  5.270 1.770 7.310 2.110 ;
        RECT  5.830 1.770 6.170 3.110 ;
        RECT  0.855 3.680 3.40 3.940 ;
        RECT  2.090 1.690 3.40 2.030 ;
        RECT  2.760 2.640 4.30 2.935 ;
        RECT  5.270 1.770 6.20 2.110 ;
    END
END ITHCX12

MACRO INX8
    CLASS CORE ;
    FOREIGN INX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.390  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.260 0.905 5.600 4.180 ;
        RECT  0.900 1.560 5.600 2.060 ;
        RECT  3.780 0.905 4.125 2.060 ;
        RECT  3.780 0.905 4.120 4.180 ;
        RECT  2.335 1.560 2.680 4.180 ;
        RECT  2.340 0.905 2.680 4.180 ;
        RECT  0.900 0.905 1.240 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.247  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.555 0.585 2.365 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.500 -0.400 4.840 1.245 ;
        RECT  3.060 -0.400 3.400 1.245 ;
        RECT  1.620 -0.400 1.960 1.245 ;
        RECT  0.180 -0.400 0.520 1.245 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.500 2.315 4.840 5.280 ;
        RECT  3.060 2.315 3.400 5.280 ;
        RECT  1.620 2.315 1.960 5.280 ;
        RECT  0.180 2.665 0.520 5.280 ;
        END
    END vdd!
END INX8

MACRO INX6
    CLASS CORE ;
    FOREIGN INX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.057  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 0.905 4.230 4.180 ;
        RECT  0.970 1.600 4.230 2.040 ;
        RECT  2.410 0.905 2.755 2.040 ;
        RECT  2.410 0.905 2.750 4.180 ;
        RECT  0.970 0.905 1.310 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.550 0.740 2.360 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.130 -0.400 3.470 1.245 ;
        RECT  1.690 -0.400 2.030 1.245 ;
        RECT  0.205 -0.400 0.550 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.130 2.270 3.470 5.280 ;
        RECT  1.690 2.270 2.030 5.280 ;
        RECT  0.210 2.660 0.550 5.280 ;
        END
    END vdd!
END INX6

MACRO INX4
    CLASS CORE ;
    FOREIGN INX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.441  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.480 0.975 2.825 4.160 ;
        RECT  1.040 1.600 2.825 2.060 ;
        RECT  1.040 0.975 1.380 4.160 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.627  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.635 0.610 2.145 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.200 -0.400 3.540 1.315 ;
        RECT  1.760 -0.400 2.100 1.315 ;
        RECT  0.320 -0.400 0.660 1.315 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.200 2.640 3.540 5.280 ;
        RECT  1.760 2.635 2.100 5.280 ;
        RECT  0.320 2.640 0.660 5.280 ;
        END
    END vdd!
END INX4

MACRO INX3
    CLASS CORE ;
    FOREIGN INX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.480 0.975 2.825 4.160 ;
        RECT  1.040 1.600 2.825 2.060 ;
        RECT  1.040 0.975 1.380 4.160 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.183  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.635 0.610 2.145 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.760 -0.400 2.100 1.315 ;
        RECT  0.320 -0.400 0.660 1.315 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.760 2.635 2.100 5.280 ;
        RECT  0.320 2.640 0.660 5.280 ;
        END
    END vdd!
END INX3

MACRO INX20
    CLASS CORE ;
    FOREIGN INX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.402  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.940 0.675 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.638  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.010 0.905 19.350 4.160 ;
        RECT  11.790 1.510 19.350 2.310 ;
        RECT  17.550 0.905 17.890 4.160 ;
        RECT  16.110 0.920 16.450 4.140 ;
        RECT  14.670 0.920 15.010 4.160 ;
        RECT  13.230 0.920 13.570 4.160 ;
        RECT  11.790 0.920 12.130 4.160 ;
        RECT  7.470 2.375 12.130 2.715 ;
        RECT  7.470 1.285 12.130 1.575 ;
        RECT  10.350 2.375 10.690 4.160 ;
        RECT  10.350 0.920 10.690 1.575 ;
        RECT  8.910 0.920 9.255 1.575 ;
        RECT  8.910 2.375 9.250 4.160 ;
        RECT  7.470 2.375 7.810 4.160 ;
        RECT  7.470 0.920 7.810 1.575 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.270 2.780 18.610 5.280 ;
        RECT  16.830 2.540 17.170 5.280 ;
        RECT  15.390 2.560 15.730 5.280 ;
        RECT  13.950 2.560 14.290 5.280 ;
        RECT  12.510 2.560 12.850 5.280 ;
        RECT  11.070 2.945 11.410 5.280 ;
        RECT  9.630 2.945 9.970 5.280 ;
        RECT  8.190 2.945 8.530 5.280 ;
        RECT  6.750 2.555 7.090 5.280 ;
        RECT  5.305 2.555 5.650 5.280 ;
        RECT  3.865 2.830 4.210 5.280 ;
        RECT  2.430 2.345 2.780 5.280 ;
        RECT  0.900 3.320 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.270 -0.400 18.610 1.245 ;
        RECT  16.830 -0.400 17.170 1.260 ;
        RECT  15.390 -0.400 15.730 1.260 ;
        RECT  13.950 -0.400 14.290 1.260 ;
        RECT  12.510 -0.400 12.850 1.260 ;
        RECT  11.070 -0.400 11.410 1.055 ;
        RECT  9.630 -0.400 9.970 1.055 ;
        RECT  8.190 -0.400 9.970 0.405 ;
        RECT  8.190 -0.400 8.530 1.055 ;
        RECT  6.750 -0.400 7.090 1.260 ;
        RECT  5.310 -0.400 5.650 1.255 ;
        RECT  3.870 -0.400 4.210 1.040 ;
        RECT  2.430 -0.400 2.775 1.245 ;
        RECT  0.895 -0.400 1.240 1.250 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.895 0.520 1.710 ;
        RECT  0.180 1.480 1.960 1.710 ;
        RECT  1.620 1.730 4.360 2.115 ;
        RECT  0.180 2.860 1.960 3.090 ;
        RECT  0.180 2.860 0.520 4.180 ;
        RECT  1.620 0.895 1.960 4.180 ;
        RECT  3.150 0.895 3.490 1.500 ;
        RECT  3.150 1.270 4.930 1.500 ;
        RECT  4.590 1.805 11.560 2.145 ;
        RECT  4.590 1.505 6.370 2.305 ;
        RECT  3.150 2.345 4.930 2.600 ;
        RECT  3.150 2.345 3.490 4.180 ;
        RECT  4.590 0.895 4.930 4.180 ;
        RECT  6.030 0.895 6.370 4.180 ;
        RECT  1.620 1.730 3.50 2.115 ;
        RECT  4.590 1.805 10.00 2.145 ;
    END
END INX20

MACRO INX2
    CLASS CORE ;
    FOREIGN INX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.003  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.775 1.030 1.135 3.160 ;
        RECT  0.755 1.030 1.135 1.410 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.851  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.030 0.545 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  1.370 3.580 1.710 5.280 ;
        RECT  0.180 3.580 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  1.370 -0.400 1.710 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
END INX2

MACRO INX16
    CLASS CORE ;
    FOREIGN INX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.878  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.880 0.920 14.220 4.160 ;
        RECT  8.135 1.490 14.220 2.190 ;
        RECT  12.440 0.920 12.785 2.190 ;
        RECT  12.440 0.920 12.780 4.160 ;
        RECT  11.000 0.920 11.340 4.160 ;
        RECT  9.560 0.920 9.905 2.190 ;
        RECT  9.560 0.920 9.900 4.160 ;
        RECT  8.120 2.390 8.460 4.160 ;
        RECT  8.135 0.920 8.460 4.160 ;
        RECT  8.120 0.920 8.460 1.580 ;
        RECT  5.240 2.390 8.460 2.730 ;
        RECT  5.240 1.285 8.460 1.580 ;
        RECT  6.680 0.920 7.025 1.580 ;
        RECT  6.680 2.390 7.020 4.160 ;
        RECT  5.240 2.390 5.580 4.160 ;
        RECT  5.240 0.920 5.580 1.580 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.767  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.625 0.690 2.050 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.600 2.840 14.955 5.280 ;
        RECT  13.160 2.440 13.500 5.280 ;
        RECT  11.720 2.440 12.060 5.280 ;
        RECT  10.280 2.440 10.620 5.280 ;
        RECT  8.840 2.440 9.180 5.280 ;
        RECT  7.400 2.960 7.740 5.280 ;
        RECT  5.960 2.960 6.300 5.280 ;
        RECT  4.515 2.390 4.860 5.280 ;
        RECT  3.075 2.830 3.420 5.280 ;
        RECT  1.640 2.900 1.990 5.280 ;
        RECT  0.200 2.900 0.540 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  14.600 -0.400 14.940 1.260 ;
        RECT  13.160 -0.400 13.500 1.260 ;
        RECT  11.720 -0.400 12.060 1.260 ;
        RECT  10.280 -0.400 10.620 1.260 ;
        RECT  8.840 -0.400 9.180 1.260 ;
        RECT  7.400 -0.400 7.740 1.055 ;
        RECT  5.960 -0.400 6.300 1.055 ;
        RECT  4.520 -0.400 4.860 1.260 ;
        RECT  3.080 -0.400 3.420 1.040 ;
        RECT  1.640 -0.400 1.985 1.245 ;
        RECT  0.195 -0.400 0.540 1.245 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.920 1.730 3.420 2.115 ;
        RECT  0.920 0.905 1.260 4.180 ;
        RECT  2.360 0.895 2.700 1.500 ;
        RECT  2.360 1.270 4.140 1.500 ;
        RECT  3.650 1.810 7.905 2.150 ;
        RECT  3.650 1.270 4.140 2.600 ;
        RECT  2.360 2.345 4.140 2.600 ;
        RECT  2.360 2.345 2.700 4.180 ;
        RECT  3.800 0.895 4.140 4.180 ;
        RECT  0.920 1.730 2.40 2.115 ;
        RECT  3.650 1.810 6.80 2.150 ;
    END
END INX16

MACRO INX12
    CLASS CORE ;
    FOREIGN INX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.815 2.035 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.690 0.905 11.030 4.180 ;
        RECT  7.530 1.480 11.030 2.080 ;
        RECT  9.210 0.905 9.555 2.080 ;
        RECT  9.210 0.905 9.550 4.180 ;
        RECT  7.770 0.905 8.110 4.180 ;
        RECT  4.850 2.360 8.110 2.650 ;
        RECT  7.530 1.270 8.110 2.650 ;
        RECT  4.850 1.270 8.110 1.560 ;
        RECT  6.290 0.905 6.635 1.560 ;
        RECT  6.290 2.360 6.630 4.180 ;
        RECT  4.850 0.905 5.195 1.560 ;
        RECT  4.850 2.360 5.190 4.180 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  11.450 -0.400 11.790 1.245 ;
        RECT  9.930 -0.400 10.270 1.245 ;
        RECT  8.490 -0.400 8.830 1.245 ;
        RECT  7.010 -0.400 7.350 1.040 ;
        RECT  5.570 -0.400 5.910 1.040 ;
        RECT  4.130 -0.400 4.470 1.245 ;
        RECT  2.690 -0.400 3.035 1.245 ;
        RECT  0.485 -0.400 0.830 1.245 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.450 2.760 11.805 5.280 ;
        RECT  9.930 2.330 10.270 5.280 ;
        RECT  8.490 2.330 8.830 5.280 ;
        RECT  7.010 2.880 7.350 5.280 ;
        RECT  5.570 2.880 5.910 5.280 ;
        RECT  4.125 2.360 4.470 5.280 ;
        RECT  2.690 2.360 3.040 5.280 ;
        RECT  0.490 2.640 0.830 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.210 1.570 1.740 2.380 ;
        RECT  1.210 0.905 1.550 4.180 ;
        RECT  1.970 1.790 7.300 2.130 ;
        RECT  1.970 0.905 2.310 4.180 ;
        RECT  3.410 0.905 3.750 4.180 ;
        RECT  1.970 1.790 6.40 2.130 ;
    END
END INX12

MACRO INX1
    CLASS CORE ;
    FOREIGN INX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.946  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.820 1.145 3.160 ;
        RECT  0.830 1.030 1.145 3.160 ;
        RECT  0.740 1.030 1.145 1.570 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.030 0.600 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        RECT  0.180 3.580 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
END INX1

MACRO INX0
    CLASS CORE ;
    FOREIGN INX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.624  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.745 2.860 1.145 3.290 ;
        RECT  0.745 1.170 1.030 3.290 ;
        RECT  0.690 1.170 1.030 1.510 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.690 0.515 2.250 ;
        RECT  0.115 1.640 0.500 2.250 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        RECT  0.180 3.980 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        RECT  0.690 -0.400 1.030 0.710 ;
        END
    END gnd!
END INX0

MACRO INCX20
    CLASS CORE ;
    FOREIGN INCX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.778  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.615 2.215 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.743  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 0.700 17.515 4.180 ;
        RECT  7.040 1.755 17.515 2.555 ;
        RECT  15.680 0.700 16.020 4.180 ;
        RECT  14.240 0.700 14.580 4.180 ;
        RECT  12.800 0.700 13.140 4.180 ;
        RECT  11.360 0.700 11.700 4.180 ;
        RECT  9.920 0.700 10.260 4.180 ;
        RECT  8.480 0.700 8.820 4.180 ;
        RECT  7.040 0.790 7.380 4.165 ;
        RECT  4.270 2.960 7.380 3.300 ;
        RECT  5.600 2.960 5.940 4.165 ;
        RECT  4.160 3.755 4.500 4.095 ;
        RECT  4.270 2.960 4.500 4.095 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.400 2.790 16.740 5.280 ;
        RECT  14.950 2.815 15.300 5.280 ;
        RECT  13.520 2.815 13.860 5.280 ;
        RECT  12.080 2.815 12.420 5.280 ;
        RECT  10.640 2.815 10.980 5.280 ;
        RECT  9.190 2.815 9.540 5.280 ;
        RECT  7.760 2.805 8.100 5.280 ;
        RECT  6.320 3.530 6.660 5.280 ;
        RECT  4.880 3.675 5.220 5.280 ;
        RECT  3.275 3.580 3.615 5.280 ;
        RECT  1.620 2.640 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.510 ;
        RECT  14.960 -0.400 15.300 1.510 ;
        RECT  13.520 -0.400 13.860 1.510 ;
        RECT  12.080 -0.400 12.420 1.510 ;
        RECT  10.640 -0.400 10.980 1.510 ;
        RECT  9.200 -0.400 9.540 1.510 ;
        RECT  7.760 -0.400 8.100 1.510 ;
        RECT  6.320 -0.400 6.660 1.170 ;
        RECT  3.250 -0.400 3.590 1.170 ;
        RECT  1.450 -0.400 1.790 0.710 ;
        RECT  0.330 -0.400 0.670 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.890 1.235 1.230 4.060 ;
        RECT  0.890 1.875 2.180 2.215 ;
        RECT  0.890 1.875 1.240 4.060 ;
        RECT  4.350 1.160 4.690 2.270 ;
        RECT  2.430 1.930 6.240 2.270 ;
        RECT  2.430 1.930 2.680 4.180 ;
        RECT  2.340 2.640 2.680 4.180 ;
        RECT  3.820 0.630 6.090 0.930 ;
        RECT  2.370 0.865 2.710 1.700 ;
        RECT  5.280 0.630 6.090 1.700 ;
        RECT  3.820 0.630 4.120 1.700 ;
        RECT  2.370 1.400 4.120 1.700 ;
        RECT  5.280 1.400 6.770 1.700 ;
        RECT  6.470 1.400 6.770 2.730 ;
        RECT  3.660 2.500 6.770 2.730 ;
        RECT  3.660 2.500 4.000 2.990 ;
        RECT  2.430 1.930 5.90 2.270 ;
        RECT  3.820 0.630 5.40 0.930 ;
        RECT  3.660 2.500 5.90 2.730 ;
    END
END INCX20

MACRO INCX16
    CLASS CORE ;
    FOREIGN INCX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.630  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.640 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.600 0.700 14.995 4.180 ;
        RECT  5.960 1.760 14.995 2.460 ;
        RECT  13.160 0.700 13.500 4.180 ;
        RECT  11.720 0.700 12.060 4.180 ;
        RECT  10.280 0.700 10.620 4.180 ;
        RECT  8.840 0.700 9.180 4.180 ;
        RECT  7.400 0.700 7.740 4.180 ;
        RECT  5.960 0.875 6.300 4.180 ;
        RECT  4.520 3.030 6.300 3.330 ;
        RECT  4.520 3.030 4.860 4.165 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.880 -0.400 14.220 1.510 ;
        RECT  12.440 -0.400 12.780 1.510 ;
        RECT  11.000 -0.400 11.340 1.510 ;
        RECT  9.560 -0.400 9.900 1.510 ;
        RECT  8.120 -0.400 8.460 1.510 ;
        RECT  6.680 -0.400 7.020 1.215 ;
        RECT  4.500 -0.400 4.840 1.070 ;
        RECT  2.540 -0.400 2.880 1.310 ;
        RECT  0.180 -0.400 0.520 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  13.880 2.740 14.220 5.280 ;
        RECT  12.430 2.690 12.780 5.280 ;
        RECT  11.000 2.690 11.340 5.280 ;
        RECT  9.560 2.690 9.900 5.280 ;
        RECT  8.120 2.690 8.460 5.280 ;
        RECT  6.670 2.690 7.020 5.280 ;
        RECT  5.240 3.560 5.580 5.280 ;
        RECT  3.065 3.825 4.140 5.280 ;
        RECT  3.065 2.760 3.405 5.280 ;
        RECT  1.620 2.640 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 0.690 1.280 2.410 ;
        RECT  0.900 2.070 2.200 2.410 ;
        RECT  0.900 0.690 1.240 3.810 ;
        RECT  1.640 0.890 1.980 1.840 ;
        RECT  1.640 1.540 2.680 1.840 ;
        RECT  2.450 1.930 5.255 2.270 ;
        RECT  2.450 1.540 2.680 3.960 ;
        RECT  2.340 2.640 2.680 3.960 ;
        RECT  3.520 0.860 3.860 1.600 ;
        RECT  5.400 0.630 5.730 1.600 ;
        RECT  3.520 1.300 5.730 1.600 ;
        RECT  5.485 0.630 5.730 2.800 ;
        RECT  3.785 2.500 5.730 2.800 ;
        RECT  3.785 2.500 4.125 3.050 ;
        RECT  2.450 1.930 4.30 2.270 ;
        RECT  3.520 1.300 4.20 1.600 ;
    END
END INCX16

MACRO INCX12
    CLASS CORE ;
    FOREIGN INCX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.956  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.220 2.135 11.590 2.420 ;
        RECT  11.250 0.700 11.590 2.420 ;
        RECT  5.490 1.820 11.590 2.420 ;
        RECT  10.730 1.820 11.070 4.180 ;
        RECT  9.810 0.700 10.150 2.420 ;
        RECT  9.290 1.820 9.630 4.180 ;
        RECT  8.315 0.700 8.710 2.420 ;
        RECT  7.850 1.820 8.190 4.180 ;
        RECT  6.930 0.700 7.270 2.420 ;
        RECT  6.410 1.820 6.750 4.180 ;
        RECT  5.490 0.700 5.830 2.420 ;
        RECT  3.470 3.180 5.460 3.460 ;
        RECT  5.220 2.135 5.460 3.460 ;
        RECT  4.970 3.180 5.310 4.180 ;
        RECT  3.470 3.180 3.810 4.120 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.580 0.760 2.020 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.530 -0.400 10.870 1.570 ;
        RECT  9.090 -0.400 9.430 1.570 ;
        RECT  7.650 -0.400 7.990 1.570 ;
        RECT  6.210 -0.400 6.550 1.570 ;
        RECT  4.240 -0.400 4.580 1.280 ;
        RECT  2.460 -0.400 2.800 1.430 ;
        RECT  0.180 -0.400 0.520 1.250 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.450 2.695 11.790 5.280 ;
        RECT  10.010 2.650 10.350 5.280 ;
        RECT  8.570 2.650 8.910 5.280 ;
        RECT  7.130 2.650 7.470 5.280 ;
        RECT  5.690 2.650 6.030 5.280 ;
        RECT  4.250 3.690 4.590 5.280 ;
        RECT  2.200 3.680 3.010 5.280 ;
        RECT  0.900 2.780 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 0.910 1.370 1.250 ;
        RECT  1.070 0.910 1.370 2.550 ;
        RECT  1.070 2.120 1.480 2.550 ;
        RECT  0.180 2.250 1.480 2.550 ;
        RECT  0.180 2.250 0.520 4.180 ;
        RECT  1.600 1.000 1.960 1.340 ;
        RECT  1.710 2.040 4.420 2.380 ;
        RECT  1.710 1.000 1.960 3.760 ;
        RECT  1.620 2.740 1.960 3.760 ;
        RECT  3.370 1.000 3.710 1.810 ;
        RECT  3.370 1.510 5.150 1.810 ;
        RECT  4.810 0.630 5.150 1.880 ;
        RECT  4.650 1.510 4.990 2.950 ;
        RECT  2.950 2.610 4.990 2.950 ;
        RECT  1.710 2.040 3.80 2.380 ;
        RECT  2.950 2.610 3.60 2.950 ;
    END
END INCX12

MACRO HAX4
    CLASS CORE ;
    FOREIGN HAX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.926  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.770 1.775 7.520 2.005 ;
        RECT  7.180 1.445 7.520 2.005 ;
        RECT  6.770 2.915 7.110 3.840 ;
        RECT  6.770 1.775 7.000 3.840 ;
        RECT  5.330 2.250 7.000 2.630 ;
        RECT  5.740 1.610 6.080 2.630 ;
        RECT  5.330 2.250 5.670 3.840 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.781  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.680 1.765 5.020 2.130 ;
        RECT  4.535 1.845 4.915 2.630 ;
        RECT  3.570 1.845 4.915 2.195 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.781  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.640 2.880 2.130 ;
        END
    END A
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.254  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.720 2.960 2.060 4.180 ;
        RECT  1.470 1.040 1.960 1.380 ;
        RECT  1.450 2.960 2.060 3.245 ;
        RECT  1.470 1.040 1.700 1.715 ;
        RECT  1.450 1.545 1.680 3.245 ;
        RECT  0.180 2.250 1.680 2.630 ;
        RECT  0.180 1.040 0.520 4.180 ;
        END
    END S
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  7.740 -0.400 8.080 0.970 ;
        RECT  6.460 -0.400 6.800 1.545 ;
        RECT  5.200 -0.400 5.540 1.250 ;
        RECT  2.340 -0.400 2.680 1.380 ;
        RECT  0.900 -0.400 1.240 1.380 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.930 2.980 9.270 5.280 ;
        RECT  7.490 2.980 7.830 5.280 ;
        RECT  6.050 2.920 6.390 5.280 ;
        RECT  4.505 3.030 4.845 5.280 ;
        RECT  2.440 2.930 2.780 5.280 ;
        RECT  0.900 3.340 1.240 5.280 ;
        RECT  0.900 2.960 1.220 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.110 1.270 4.100 1.615 ;
        RECT  3.110 1.270 3.340 2.810 ;
        RECT  1.910 2.360 3.340 2.700 ;
        RECT  3.110 2.550 3.930 2.810 ;
        RECT  3.590 2.550 3.930 3.880 ;
        RECT  3.060 0.700 4.820 1.040 ;
        RECT  4.480 0.700 4.820 1.535 ;
        RECT  8.930 0.700 9.270 2.575 ;
        RECT  7.250 2.235 9.270 2.575 ;
        RECT  8.210 2.235 8.550 3.840 ;
        RECT  7.250 2.235 8.30 2.575 ;
    END
END HAX4

MACRO HAX2
    CLASS CORE ;
    FOREIGN HAX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALAREA 0.474  LAYER MET1  ;
        ANTENNAGATEAREA 0.745  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.170 3.520 6.805 4.100 ;
        RECT  4.000 1.765 4.340 2.075 ;
        RECT  2.850 1.845 4.335 2.130 ;
        RECT  2.850 1.845 3.190 2.195 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.903  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.100 1.445 5.630 1.785 ;
        RECT  4.955 1.755 5.330 1.970 ;
        RECT  4.880 2.570 5.220 3.840 ;
        RECT  4.535 2.250 5.185 2.630 ;
        RECT  4.955 1.755 5.185 3.840 ;
        END
    END CO
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.745  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.640 2.160 2.130 ;
        END
    END A
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 2.960 1.240 3.880 ;
        RECT  0.750 1.105 1.240 1.445 ;
        RECT  0.750 1.105 0.980 3.245 ;
        RECT  0.125 2.250 0.980 2.630 ;
        END
    END S
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.850 -0.400 6.190 0.970 ;
        RECT  4.520 -0.400 4.860 1.545 ;
        RECT  1.660 -0.400 2.000 1.410 ;
        RECT  0.180 -0.400 0.520 1.425 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 3.080 7.380 5.280 ;
        RECT  5.600 3.100 5.940 5.280 ;
        RECT  3.550 3.030 4.500 5.280 ;
        RECT  1.620 3.000 1.960 5.280 ;
        RECT  0.180 2.960 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.390 1.270 3.420 1.615 ;
        RECT  2.390 1.270 2.620 2.810 ;
        RECT  1.210 2.390 2.620 2.730 ;
        RECT  2.390 2.550 3.110 2.810 ;
        RECT  2.770 2.550 3.110 3.880 ;
        RECT  2.380 0.700 4.140 1.040 ;
        RECT  3.800 0.700 4.140 1.510 ;
        RECT  5.445 2.170 7.380 2.415 ;
        RECT  7.040 0.700 7.380 2.415 ;
        RECT  5.415 2.185 7.380 2.415 ;
        RECT  5.445 2.170 6.660 2.470 ;
        RECT  6.320 2.170 6.660 3.290 ;
    END
END HAX2

MACRO HAX1
    CLASS CORE ;
    FOREIGN HAX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.710 1.610 4.370 1.950 ;
        RECT  3.620 2.250 3.960 3.880 ;
        RECT  3.710 1.610 3.960 3.880 ;
        RECT  3.200 2.250 3.960 2.630 ;
        END
    END CO
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.677  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 1.675 1.890 2.145 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.695  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.910 3.520 5.545 4.100 ;
        END
    END B
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.757  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.240 1.360 1.080 1.700 ;
        RECT  0.330 2.850 0.670 3.770 ;
        RECT  0.240 1.360 0.505 3.135 ;
        RECT  0.125 2.250 0.505 2.630 ;
        END
    END S
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 3.080 6.120 5.280 ;
        RECT  4.340 3.100 4.680 5.280 ;
        RECT  2.920 2.960 3.260 5.280 ;
        RECT  1.050 2.890 1.390 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.590 -0.400 4.930 0.970 ;
        RECT  2.000 -0.400 2.340 0.985 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.280 0.700 1.620 1.040 ;
        RECT  1.310 0.700 1.620 1.445 ;
        RECT  1.310 1.215 3.020 1.445 ;
        RECT  2.680 1.215 3.020 1.560 ;
        RECT  3.250 1.000 3.750 1.340 ;
        RECT  3.250 1.000 3.480 2.020 ;
        RECT  2.310 1.790 3.480 2.020 ;
        RECT  0.810 2.320 1.150 2.660 ;
        RECT  0.810 2.375 2.540 2.660 ;
        RECT  2.310 1.790 2.540 3.310 ;
        RECT  2.200 2.375 2.540 3.310 ;
        RECT  5.780 0.700 6.120 2.415 ;
        RECT  4.270 2.180 6.120 2.415 ;
        RECT  4.270 2.180 5.400 2.470 ;
        RECT  5.060 2.180 5.400 3.290 ;
    END
END HAX1

MACRO HAX0
    CLASS CORE ;
    FOREIGN HAX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.570 1.370 4.215 1.660 ;
        RECT  3.570 1.370 3.800 2.580 ;
        RECT  3.385 2.250 3.725 3.060 ;
        RECT  3.275 2.250 3.725 2.630 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.845 3.470 2.395 3.920 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.288  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.315 0.630 5.765 0.915 ;
        RECT  5.165 1.030 5.545 1.410 ;
        RECT  5.315 0.630 5.545 1.410 ;
        END
    END A
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.240 2.640 0.635 2.980 ;
        RECT  0.185 1.170 0.525 1.510 ;
        RECT  0.240 1.170 0.505 2.980 ;
        RECT  0.125 2.250 0.505 2.630 ;
        RECT  0.185 1.170 0.505 2.630 ;
        END
    END S
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.585 2.860 5.925 5.280 ;
        RECT  3.985 3.510 4.325 5.280 ;
        RECT  2.685 3.380 3.025 5.280 ;
        RECT  0.295 3.415 1.435 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.475 -0.400 4.815 0.970 ;
        RECT  1.825 -0.400 2.165 0.915 ;
        RECT  0.185 -0.400 0.525 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.025 0.980 1.365 1.375 ;
        RECT  2.585 0.960 2.880 1.375 ;
        RECT  1.025 1.145 2.880 1.375 ;
        RECT  3.110 0.670 3.735 1.010 ;
        RECT  3.110 0.670 3.340 1.835 ;
        RECT  0.735 1.605 3.340 1.835 ;
        RECT  0.735 1.605 1.045 1.945 ;
        RECT  2.085 1.605 2.425 2.980 ;
        RECT  5.775 1.170 6.060 2.120 ;
        RECT  4.030 1.890 6.060 2.120 ;
        RECT  4.030 1.890 4.315 2.230 ;
        RECT  4.785 1.890 5.125 3.210 ;
        RECT  0.735 1.605 2.20 1.835 ;
        RECT  4.030 1.890 5.50 2.120 ;
    END
END HAX0

MACRO FEEDCAP7LP
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP7LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.275 -0.400 3.615 1.310 ;
        RECT  0.795 -0.400 1.135 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.255 4.190 3.135 5.280 ;
        END
    END vdd!
END FEEDCAP7LP

MACRO FEEDCAP7
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.890 -0.400 4.230 0.710 ;
        RECT  0.165 -0.400 0.520 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  0.975 4.190 3.490 5.280 ;
        END
    END vdd!
END FEEDCAP7

MACRO FEEDCAP5LP
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP5LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.015 -0.400 2.355 1.310 ;
        RECT  0.795 -0.400 1.135 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.640 4.190 2.530 5.280 ;
        END
    END vdd!
END FEEDCAP5LP

MACRO FEEDCAP5
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP5 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 0.710 ;
        RECT  0.165 -0.400 1.025 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.125 4.170 2.985 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
END FEEDCAP5

MACRO FEEDCAP3
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  0.140 -0.400 1.750 1.060 ;
        RECT  0.140 -0.400 0.520 2.700 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  0.180 3.840 1.745 5.280 ;
        RECT  1.380 1.895 1.745 5.280 ;
        END
    END vdd!
END FEEDCAP3

MACRO FEEDCAP25LP
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP25LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  14.615 -0.400 14.955 1.310 ;
        RECT  12.115 -0.400 12.455 1.310 ;
        RECT  8.335 -0.400 8.675 1.310 ;
        RECT  4.555 -0.400 4.895 1.310 ;
        RECT  0.795 -0.400 1.135 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  1.380 4.190 14.455 5.280 ;
        END
    END vdd!
END FEEDCAP25LP

MACRO FEEDCAP25
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP25 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.230 -0.400 15.570 0.710 ;
        RECT  11.200 -0.400 11.560 0.715 ;
        RECT  7.695 -0.400 8.055 0.710 ;
        RECT  4.190 -0.400 4.550 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  1.305 4.190 14.490 5.280 ;
        END
    END vdd!
END FEEDCAP25

MACRO FEEDCAP2
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        RECT  0.140 -0.400 1.120 1.060 ;
        RECT  0.140 -0.400 0.520 2.700 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        RECT  0.180 3.840 1.115 5.280 ;
        RECT  0.750 1.895 1.115 5.280 ;
        END
    END vdd!
END FEEDCAP2

MACRO FEEDCAP15LP
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP15LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.315 -0.400 8.655 1.310 ;
        RECT  4.555 -0.400 4.895 1.310 ;
        RECT  0.795 -0.400 1.135 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  1.310 4.190 8.205 5.280 ;
        END
    END vdd!
END FEEDCAP15LP

MACRO FEEDCAP15
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP15 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.930 -0.400 9.270 0.710 ;
        RECT  4.545 -0.400 4.905 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  1.305 4.190 8.190 5.280 ;
        END
    END vdd!
END FEEDCAP15

MACRO FEEDCAP10LP
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP10LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.165 -0.400 5.505 1.310 ;
        RECT  0.795 -0.400 1.135 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  1.195 4.190 5.125 5.280 ;
        END
    END vdd!
END FEEDCAP10LP

MACRO FEEDCAP10
    CLASS CORE SPACER ;
    FOREIGN FEEDCAP10 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  1.495 4.190 4.850 5.280 ;
        END
    END vdd!
END FEEDCAP10

MACRO FEED7
    CLASS CORE SPACER ;
    FOREIGN FEED7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        END
    END gnd!
END FEED7

MACRO FEED5
    CLASS CORE SPACER ;
    FOREIGN FEED5 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        END
    END gnd!
END FEED5

MACRO FEED3
    CLASS CORE SPACER ;
    FOREIGN FEED3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        END
    END gnd!
END FEED3

MACRO FEED25
    CLASS CORE SPACER ;
    FOREIGN FEED25 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        END
    END gnd!
END FEED25

MACRO FEED2
    CLASS CORE SPACER ;
    FOREIGN FEED2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        END
    END gnd!
END FEED2

MACRO FEED15
    CLASS CORE SPACER ;
    FOREIGN FEED15 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        END
    END gnd!
END FEED15

MACRO FEED10
    CLASS CORE SPACER ;
    FOREIGN FEED10 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        END
    END gnd!
END FEED10

MACRO FEED1
    CLASS CORE SPACER ;
    FOREIGN FEED1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.630 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 0.630 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 0.630 0.400 ;
        END
    END gnd!
END FEED1

MACRO FAX4
    CLASS CORE ;
    FOREIGN FAX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 0.700 1.960 4.180 ;
        RECT  1.385 2.250 1.960 2.630 ;
        RECT  0.180 2.250 1.960 2.480 ;
        RECT  0.180 0.700 0.520 4.180 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.023  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.415 1.130 10.905 1.470 ;
        RECT  10.415 1.130 10.645 1.690 ;
        RECT  8.595 2.570 10.610 2.855 ;
        RECT  10.205 2.250 10.610 2.855 ;
        RECT  10.380 1.565 10.610 2.855 ;
        RECT  9.125 1.110 9.465 2.855 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.123  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.840 2.610 12.710 2.895 ;
        RECT  12.095 2.555 12.710 2.895 ;
        RECT  12.095 2.240 12.475 2.895 ;
        RECT  8.135 3.085 11.070 3.315 ;
        RECT  10.840 2.610 11.070 3.315 ;
        RECT  7.260 3.080 8.365 3.310 ;
        RECT  6.175 3.210 7.490 3.440 ;
        RECT  6.175 2.135 7.140 2.385 ;
        RECT  6.175 2.135 6.405 3.440 ;
        RECT  3.225 2.540 6.405 2.825 ;
        RECT  3.225 2.540 3.565 2.855 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.454  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.690 4.015 14.365 4.250 ;
        RECT  13.985 3.470 14.365 4.250 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.540 2.045 14.995 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  14.600 2.875 14.940 5.280 ;
        RECT  12.030 3.705 12.370 5.280 ;
        RECT  10.590 3.545 10.930 5.280 ;
        RECT  9.260 3.545 9.600 5.280 ;
        RECT  5.145 3.540 5.485 5.280 ;
        RECT  3.705 3.575 4.045 5.280 ;
        RECT  2.340 3.760 2.680 5.280 ;
        RECT  0.900 2.900 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  13.880 -0.400 14.220 1.340 ;
        RECT  11.290 -0.400 11.630 1.470 ;
        RECT  9.845 -0.400 10.185 1.440 ;
        RECT  8.405 -0.400 8.745 1.450 ;
        RECT  5.900 -0.400 6.240 0.985 ;
        RECT  4.465 -0.400 4.805 1.495 ;
        RECT  2.340 -0.400 2.680 1.100 ;
        RECT  0.900 -0.400 1.240 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  5.180 0.700 5.520 1.445 ;
        RECT  6.830 1.160 7.170 1.445 ;
        RECT  5.180 1.215 7.170 1.445 ;
        RECT  2.880 1.460 3.220 2.110 ;
        RECT  5.235 1.675 8.000 1.905 ;
        RECT  7.660 1.155 8.000 1.905 ;
        RECT  2.360 1.880 5.465 2.110 ;
        RECT  2.360 1.880 2.700 2.220 ;
        RECT  7.370 1.675 7.600 2.845 ;
        RECT  6.745 2.615 7.600 2.845 ;
        RECT  6.745 2.615 7.060 2.965 ;
        RECT  6.745 2.615 7.030 2.980 ;
        RECT  4.425 3.060 5.945 3.310 ;
        RECT  2.985 3.115 4.765 3.345 ;
        RECT  2.985 3.085 3.325 3.400 ;
        RECT  5.715 3.060 5.945 3.900 ;
        RECT  4.425 3.060 4.765 3.870 ;
        RECT  7.710 3.540 8.005 3.900 ;
        RECT  5.715 3.670 8.005 3.900 ;
        RECT  11.310 3.135 13.070 3.475 ;
        RECT  11.310 3.135 11.650 3.585 ;
        RECT  12.440 1.130 12.780 2.010 ;
        RECT  10.860 1.775 12.780 2.010 ;
        RECT  10.860 1.780 13.170 2.010 ;
        RECT  10.840 1.815 11.700 2.045 ;
        RECT  10.840 1.815 11.180 2.100 ;
        RECT  12.940 1.780 13.170 2.470 ;
        RECT  12.940 2.240 13.790 2.470 ;
        RECT  13.450 2.240 13.790 3.045 ;
        RECT  13.450 2.240 13.755 3.785 ;
        RECT  13.160 1.265 13.630 1.550 ;
        RECT  13.400 1.265 13.630 1.800 ;
        RECT  14.600 1.050 14.940 1.800 ;
        RECT  13.400 1.570 14.940 1.800 ;
        RECT  5.235 1.675 7.00 1.905 ;
        RECT  2.360 1.880 4.40 2.110 ;
        RECT  5.715 3.670 7.60 3.900 ;
        RECT  10.860 1.780 12.50 2.010 ;
    END
END FAX4

MACRO FAX2
    CLASS CORE ;
    FOREIGN FAX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.454  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.800 4.015 12.475 4.250 ;
        RECT  12.095 3.470 12.475 4.250 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.472  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.650 2.045 13.105 2.630 ;
        END
    END A
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.123  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 2.240 11.090 2.475 ;
        RECT  9.015 2.510 10.585 2.740 ;
        RECT  10.205 2.240 10.585 2.740 ;
        RECT  7.355 3.105 9.245 3.335 ;
        RECT  9.015 2.510 9.245 3.335 ;
        RECT  6.435 3.075 7.585 3.305 ;
        RECT  5.515 3.440 6.665 3.670 ;
        RECT  6.435 3.075 6.665 3.670 ;
        RECT  5.515 2.135 6.315 2.385 ;
        RECT  5.515 2.135 5.745 3.670 ;
        RECT  2.400 2.540 5.745 2.825 ;
        RECT  2.400 2.540 2.740 2.855 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.395 1.130 8.925 1.470 ;
        RECT  8.100 2.590 8.695 2.875 ;
        RECT  8.315 2.255 8.695 2.875 ;
        RECT  8.315 2.250 8.625 2.875 ;
        RECT  8.395 1.130 8.625 2.875 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 3.260 1.240 4.170 ;
        RECT  0.900 0.820 1.240 1.160 ;
        RECT  0.900 0.820 1.185 4.170 ;
        RECT  0.755 2.250 1.185 2.630 ;
        END
    END S
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.990 -0.400 12.330 1.160 ;
        RECT  9.335 -0.400 9.675 1.470 ;
        RECT  7.825 -0.400 8.165 1.450 ;
        RECT  5.075 -0.400 5.415 0.985 ;
        RECT  3.640 -0.400 3.980 1.495 ;
        RECT  1.660 -0.400 2.000 0.710 ;
        RECT  0.180 -0.400 0.520 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  12.710 2.875 13.050 5.280 ;
        RECT  10.140 3.430 10.480 5.280 ;
        RECT  8.660 3.910 9.000 5.280 ;
        RECT  7.540 3.910 7.880 5.280 ;
        RECT  4.320 3.540 4.660 5.280 ;
        RECT  2.880 3.575 3.220 5.280 ;
        RECT  1.620 3.760 1.960 5.280 ;
        RECT  0.180 3.260 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  4.355 0.700 4.695 1.445 ;
        RECT  6.005 1.105 6.345 1.445 ;
        RECT  4.355 1.215 6.345 1.445 ;
        RECT  1.990 1.590 2.330 2.110 ;
        RECT  1.415 1.675 2.330 2.110 ;
        RECT  4.830 1.675 7.175 1.905 ;
        RECT  6.835 1.155 7.175 1.905 ;
        RECT  1.415 1.880 5.060 2.110 ;
        RECT  6.700 1.675 6.930 2.845 ;
        RECT  5.975 2.615 6.930 2.845 ;
        RECT  5.975 2.615 6.205 3.210 ;
        RECT  3.600 3.060 5.120 3.310 ;
        RECT  2.160 3.115 3.940 3.345 ;
        RECT  2.160 3.085 2.500 3.400 ;
        RECT  3.600 3.060 3.940 3.870 ;
        RECT  4.890 3.060 5.120 4.130 ;
        RECT  6.895 3.535 7.180 4.130 ;
        RECT  4.890 3.900 7.180 4.130 ;
        RECT  9.475 2.970 11.180 3.200 ;
        RECT  10.840 2.705 11.180 3.785 ;
        RECT  9.475 2.970 9.760 3.880 ;
        RECT  9.420 3.540 9.760 3.880 ;
        RECT  10.510 1.130 10.850 2.010 ;
        RECT  8.855 1.760 10.850 2.010 ;
        RECT  8.855 1.780 11.480 2.010 ;
        RECT  8.855 1.760 9.810 2.045 ;
        RECT  11.310 1.850 11.900 2.080 ;
        RECT  8.860 1.760 9.195 2.090 ;
        RECT  11.615 1.850 11.900 3.215 ;
        RECT  11.560 2.875 11.845 3.785 ;
        RECT  11.560 3.445 11.865 3.785 ;
        RECT  11.230 1.265 11.570 1.550 ;
        RECT  11.230 1.320 11.820 1.550 ;
        RECT  12.710 1.050 13.050 1.620 ;
        RECT  11.650 1.390 13.050 1.620 ;
        RECT  4.830 1.675 6.10 1.905 ;
        RECT  1.415 1.880 4.40 2.110 ;
        RECT  4.890 3.900 6.60 4.130 ;
        RECT  8.855 1.780 10.40 2.010 ;
    END
END FAX2

MACRO FAX1
    CLASS CORE ;
    FOREIGN FAX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.931  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.700 2.400 10.030 2.645 ;
        RECT  8.945 2.250 9.325 2.645 ;
        RECT  4.970 3.225 7.930 3.455 ;
        RECT  7.700 2.400 7.930 3.455 ;
        RECT  5.080 2.245 5.530 2.505 ;
        RECT  4.970 2.255 5.200 3.455 ;
        RECT  1.930 2.255 5.200 2.540 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.228  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.390 2.045 11.845 2.630 ;
        END
    END A
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.610 3.850 ;
        RECT  0.270 2.720 0.610 3.850 ;
        RECT  0.270 1.230 0.610 1.570 ;
        RECT  0.270 1.230 0.555 3.850 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.228  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.540 4.015 11.215 4.250 ;
        RECT  10.835 3.470 11.215 4.250 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.725  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 0.995 7.655 1.470 ;
        RECT  6.840 2.710 7.180 2.995 ;
        RECT  6.950 0.995 7.180 2.995 ;
        END
    END CO
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.690 -0.400 11.030 1.215 ;
        RECT  8.035 -0.400 8.375 1.470 ;
        RECT  4.790 -0.400 5.130 1.095 ;
        RECT  3.270 -0.400 3.610 1.340 ;
        RECT  0.990 -0.400 1.330 1.565 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.450 2.875 11.790 5.280 ;
        RECT  8.880 3.430 9.220 5.280 ;
        RECT  7.400 3.910 7.740 5.280 ;
        RECT  3.850 3.360 4.190 5.280 ;
        RECT  2.410 3.360 2.750 5.280 ;
        RECT  0.990 2.720 1.330 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.990 0.930 4.330 1.555 ;
        RECT  5.550 1.110 5.835 1.555 ;
        RECT  3.990 1.325 5.835 1.555 ;
        RECT  1.690 2.845 4.740 3.130 ;
        RECT  4.510 2.845 4.740 3.970 ;
        RECT  1.690 2.845 2.030 3.700 ;
        RECT  3.130 2.845 3.470 3.700 ;
        RECT  4.510 3.685 6.570 3.970 ;
        RECT  6.065 1.110 6.610 1.450 ;
        RECT  1.690 1.160 2.030 2.015 ;
        RECT  1.690 1.785 6.295 2.015 ;
        RECT  6.065 1.110 6.295 2.015 ;
        RECT  0.785 1.795 1.975 2.025 ;
        RECT  0.785 1.795 1.090 2.210 ;
        RECT  5.760 1.785 5.990 2.995 ;
        RECT  5.430 2.735 5.990 2.995 ;
        RECT  8.160 2.970 9.920 3.200 ;
        RECT  9.580 2.875 9.920 3.785 ;
        RECT  8.160 2.970 8.545 3.880 ;
        RECT  9.210 1.130 9.550 2.020 ;
        RECT  7.410 1.760 9.550 2.020 ;
        RECT  7.410 1.790 9.785 2.020 ;
        RECT  7.410 1.760 8.775 2.045 ;
        RECT  7.410 1.760 7.750 2.100 ;
        RECT  9.555 1.940 10.640 2.170 ;
        RECT  10.300 1.940 10.640 3.215 ;
        RECT  10.300 1.940 10.585 3.785 ;
        RECT  10.300 3.445 10.605 3.785 ;
        RECT  9.930 1.130 10.270 1.470 ;
        RECT  11.450 1.130 11.790 1.675 ;
        RECT  9.985 1.445 11.790 1.675 ;
        RECT  1.690 2.845 3.80 3.130 ;
        RECT  4.510 3.685 5.40 3.970 ;
        RECT  1.690 1.785 5.40 2.015 ;
        RECT  7.410 1.760 8.30 2.020 ;
        RECT  7.410 1.790 8.20 2.020 ;
    END
END FAX1

MACRO FAX0
    CLASS CORE ;
    FOREIGN FAX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.120 1.330 6.945 1.560 ;
        RECT  6.575 1.265 6.945 1.560 ;
        RECT  5.795 2.860 6.350 3.275 ;
        RECT  6.120 1.330 6.350 3.275 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.775 2.110 10.585 2.630 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.436  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.780 2.400 9.085 2.630 ;
        RECT  7.685 2.250 9.085 2.630 ;
        RECT  4.175 3.505 7.010 3.735 ;
        RECT  6.780 2.400 7.010 3.735 ;
        RECT  4.175 2.410 4.695 2.750 ;
        RECT  4.175 2.105 4.405 3.735 ;
        RECT  1.365 2.105 4.405 2.445 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.572  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.705 1.030 9.325 1.410 ;
        RECT  8.705 0.650 9.045 1.410 ;
        END
    END A
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.240 2.850 0.635 3.190 ;
        RECT  0.185 1.170 0.525 1.510 ;
        RECT  0.240 1.170 0.505 3.190 ;
        RECT  0.125 2.250 0.505 2.630 ;
        RECT  0.185 1.170 0.505 2.630 ;
        END
    END S
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.145 3.850 10.485 5.280 ;
        RECT  8.015 3.805 8.355 5.280 ;
        RECT  6.495 3.965 6.835 5.280 ;
        RECT  2.985 3.450 3.315 5.280 ;
        RECT  1.655 3.430 1.995 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.915 -0.400 10.255 1.695 ;
        RECT  9.275 -0.400 10.255 0.710 ;
        RECT  7.165 -0.400 7.535 0.970 ;
        RECT  4.345 -0.400 4.685 0.915 ;
        RECT  2.745 -0.400 3.085 1.340 ;
        RECT  0.185 -0.400 0.525 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.545 0.740 3.885 1.375 ;
        RECT  5.145 0.800 5.430 1.375 ;
        RECT  3.545 1.145 5.430 1.375 ;
        RECT  1.095 2.695 3.945 3.035 ;
        RECT  3.715 2.695 3.945 4.250 ;
        RECT  3.715 3.965 5.550 4.250 ;
        RECT  5.660 0.630 6.295 0.970 ;
        RECT  1.030 1.150 1.350 1.835 ;
        RECT  5.660 0.630 5.890 1.835 ;
        RECT  0.735 1.605 5.890 1.835 ;
        RECT  0.735 1.605 1.035 2.430 ;
        RECT  5.130 1.605 5.360 3.275 ;
        RECT  4.635 2.990 5.360 3.275 ;
        RECT  7.255 3.095 8.855 3.435 ;
        RECT  7.255 3.095 7.595 3.875 ;
        RECT  8.410 1.640 8.750 2.020 ;
        RECT  6.580 1.790 9.545 2.020 ;
        RECT  6.580 1.790 6.920 2.170 ;
        RECT  9.315 1.790 9.545 4.190 ;
        RECT  9.075 3.850 9.545 4.190 ;
        RECT  1.095 2.695 2.80 3.035 ;
        RECT  0.735 1.605 4.80 1.835 ;
        RECT  6.580 1.790 8.80 2.020 ;
    END
END FAX0

MACRO EO3X4
    CLASS CORE ;
    FOREIGN EO3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.922  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.660 2.920 11.160 3.260 ;
        RECT  9.550 1.365 11.160 1.715 ;
        RECT  10.820 1.355 11.160 1.715 ;
        RECT  10.205 1.365 10.585 3.260 ;
        RECT  9.550 1.360 9.890 1.715 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.565  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.375 3.240 ;
        RECT  4.035 2.420 4.375 3.240 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 2.675 3.000 ;
        RECT  2.015 2.250 2.675 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.240 3.560 10.580 5.280 ;
        RECT  9.005 3.555 9.345 5.280 ;
        RECT  6.230 3.370 6.570 5.280 ;
        RECT  4.725 3.760 5.065 5.280 ;
        RECT  2.200 3.840 2.545 5.280 ;
        RECT  0.510 3.960 0.850 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.185 -0.400 10.525 1.135 ;
        RECT  8.950 -0.400 9.290 1.085 ;
        RECT  7.670 -0.400 8.010 1.340 ;
        RECT  5.760 -0.400 6.100 1.510 ;
        RECT  3.575 -0.400 3.955 1.040 ;
        RECT  1.630 -0.400 1.970 1.340 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.485 3.380 3.215 3.610 ;
        RECT  2.935 3.380 3.215 4.180 ;
        RECT  2.935 3.840 3.260 4.180 ;
        RECT  1.485 3.380 1.825 4.185 ;
        RECT  0.905 1.790 3.345 2.020 ;
        RECT  3.000 1.790 3.345 2.130 ;
        RECT  0.905 1.000 1.235 2.985 ;
        RECT  4.185 0.630 5.390 0.940 ;
        RECT  2.805 1.000 3.160 1.560 ;
        RECT  4.185 0.630 4.465 1.560 ;
        RECT  2.805 1.270 4.465 1.560 ;
        RECT  3.575 1.270 3.805 2.595 ;
        RECT  3.445 2.365 3.675 3.700 ;
        RECT  3.635 3.470 3.985 4.040 ;
        RECT  5.500 2.910 7.305 3.140 ;
        RECT  5.500 2.910 5.865 4.180 ;
        RECT  6.940 2.910 7.305 4.180 ;
        RECT  4.735 1.170 5.075 2.950 ;
        RECT  4.735 2.300 7.440 2.640 ;
        RECT  4.735 2.300 5.090 2.950 ;
        RECT  6.950 1.270 7.290 1.800 ;
        RECT  6.950 1.570 8.020 1.800 ;
        RECT  7.670 1.570 8.020 2.290 ;
        RECT  7.670 1.950 8.200 2.290 ;
        RECT  7.670 1.570 8.010 4.180 ;
        RECT  8.370 1.360 8.725 1.700 ;
        RECT  8.430 1.945 9.650 2.285 ;
        RECT  8.430 1.360 8.725 3.260 ;
        RECT  8.370 2.915 8.725 3.260 ;
        RECT  0.905 1.790 2.30 2.020 ;
        RECT  4.735 2.300 6.70 2.640 ;
    END
END EO3X4

MACRO EO3X2
    CLASS CORE ;
    FOREIGN EO3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.750 9.970 3.560 ;
        RECT  9.740 1.250 9.970 3.560 ;
        RECT  9.630 1.250 9.970 1.590 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.375 3.240 ;
        RECT  4.035 2.420 4.375 3.240 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 2.675 3.000 ;
        RECT  2.015 2.250 2.675 2.630 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 0.720 ;
        RECT  9.065 -0.400 9.410 0.720 ;
        RECT  7.610 -0.400 7.950 1.510 ;
        RECT  5.620 -0.400 5.960 1.510 ;
        RECT  3.575 -0.400 3.955 1.040 ;
        RECT  1.630 -0.400 1.970 1.340 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 3.960 10.530 5.280 ;
        RECT  9.070 3.960 9.410 5.280 ;
        RECT  6.230 3.660 6.570 5.280 ;
        RECT  4.725 3.760 5.065 5.280 ;
        RECT  2.200 3.840 2.545 5.280 ;
        RECT  0.510 3.960 0.850 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.485 3.380 3.215 3.610 ;
        RECT  2.935 3.380 3.215 4.180 ;
        RECT  2.935 3.840 3.260 4.180 ;
        RECT  1.485 3.380 1.825 4.185 ;
        RECT  0.905 1.790 3.345 2.020 ;
        RECT  3.000 1.790 3.345 2.130 ;
        RECT  0.905 1.000 1.235 2.985 ;
        RECT  4.185 0.630 5.390 0.940 ;
        RECT  2.805 1.000 3.160 1.560 ;
        RECT  4.185 0.630 4.465 1.560 ;
        RECT  2.805 1.270 4.465 1.560 ;
        RECT  3.575 1.270 3.805 2.595 ;
        RECT  3.445 2.365 3.675 3.700 ;
        RECT  3.635 3.470 3.985 4.040 ;
        RECT  5.500 3.190 7.305 3.420 ;
        RECT  5.500 3.190 5.865 4.005 ;
        RECT  6.940 3.190 7.305 4.005 ;
        RECT  4.735 1.170 5.075 2.950 ;
        RECT  4.735 2.405 7.480 2.745 ;
        RECT  4.735 2.405 5.090 2.950 ;
        RECT  6.810 1.170 7.150 2.175 ;
        RECT  6.810 1.945 8.150 2.175 ;
        RECT  7.710 1.945 8.150 2.285 ;
        RECT  7.710 1.945 8.010 4.150 ;
        RECT  7.670 3.800 8.010 4.150 ;
        RECT  8.310 1.250 8.695 1.590 ;
        RECT  8.380 1.945 9.510 2.285 ;
        RECT  8.380 1.250 8.695 3.560 ;
        RECT  8.310 2.640 8.695 3.560 ;
        RECT  0.905 1.790 2.30 2.020 ;
        RECT  4.735 2.405 6.70 2.745 ;
    END
END EO3X2

MACRO EO3X1
    CLASS CORE ;
    FOREIGN EO3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.093  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 2.820 8.065 4.180 ;
        RECT  7.725 1.570 8.065 4.180 ;
        RECT  7.685 1.570 8.065 2.020 ;
        RECT  6.950 1.570 8.065 1.800 ;
        RECT  6.950 1.195 7.290 1.800 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.565  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.375 3.240 ;
        RECT  4.035 2.420 4.375 3.240 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 2.675 3.000 ;
        RECT  2.015 2.250 2.675 2.630 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 1.340 ;
        RECT  5.800 -0.400 6.140 1.520 ;
        RECT  3.575 -0.400 3.955 1.040 ;
        RECT  1.630 -0.400 1.970 1.340 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.230 3.370 6.570 5.280 ;
        RECT  4.725 3.760 5.065 5.280 ;
        RECT  2.200 3.840 2.545 5.280 ;
        RECT  0.510 3.960 0.850 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.485 3.380 3.215 3.610 ;
        RECT  2.935 3.380 3.215 4.180 ;
        RECT  2.935 3.840 3.260 4.180 ;
        RECT  1.485 3.380 1.825 4.185 ;
        RECT  0.905 1.790 3.345 2.020 ;
        RECT  3.000 1.790 3.345 2.130 ;
        RECT  0.905 1.000 1.235 2.985 ;
        RECT  4.185 0.630 5.390 0.940 ;
        RECT  2.805 1.000 3.160 1.560 ;
        RECT  4.185 0.630 4.465 1.560 ;
        RECT  2.805 1.270 4.465 1.560 ;
        RECT  3.575 1.270 3.805 2.595 ;
        RECT  3.445 2.365 3.675 3.700 ;
        RECT  3.635 3.470 3.985 4.040 ;
        RECT  5.500 2.910 7.305 3.140 ;
        RECT  5.500 2.910 5.865 4.180 ;
        RECT  6.940 2.910 7.305 4.180 ;
        RECT  4.735 1.170 5.075 2.950 ;
        RECT  4.735 2.300 7.475 2.640 ;
        RECT  4.735 2.300 5.090 2.950 ;
        RECT  0.905 1.790 2.10 2.020 ;
        RECT  4.735 2.300 6.30 2.640 ;
    END
END EO3X1

MACRO EO3X0
    CLASS CORE ;
    FOREIGN EO3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 2.090 3.705 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.604  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.935 2.850 5.545 3.190 ;
        RECT  5.165 1.170 5.545 3.190 ;
        RECT  4.770 1.170 5.545 1.510 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.209  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.755 2.250 2.395 2.635 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.209  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.635 3.025 2.210 ;
        RECT  2.600 1.635 3.025 2.145 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.270 4.110 4.610 5.280 ;
        RECT  2.710 2.860 3.050 5.280 ;
        RECT  1.110 3.835 1.450 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.300 -0.400 5.110 0.710 ;
        RECT  2.700 -0.400 3.040 1.405 ;
        RECT  0.630 -0.400 1.440 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.970 1.510 ;
        RECT  0.180 1.170 0.520 4.250 ;
        RECT  0.780 2.850 1.065 3.605 ;
        RECT  0.780 3.375 2.250 3.605 ;
        RECT  1.910 3.375 2.250 4.080 ;
        RECT  1.900 0.630 2.250 1.305 ;
        RECT  1.295 1.075 2.250 1.305 ;
        RECT  0.750 2.160 1.525 2.500 ;
        RECT  1.295 1.075 1.525 3.145 ;
        RECT  1.295 2.865 1.820 3.145 ;
        RECT  3.490 0.630 3.840 1.305 ;
        RECT  3.490 1.075 4.415 1.305 ;
        RECT  4.080 1.075 4.415 3.190 ;
        RECT  4.080 2.160 4.935 2.500 ;
        RECT  4.080 2.160 4.420 3.190 ;
        RECT  3.510 3.570 5.285 3.880 ;
        RECT  4.945 3.570 5.285 3.910 ;
        RECT  3.510 3.570 3.850 4.120 ;
    END
END EO3X0

MACRO EO2X4
    CLASS CORE ;
    FOREIGN EO2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.922  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.880 2.920 7.380 3.260 ;
        RECT  5.770 1.365 7.380 1.715 ;
        RECT  7.040 1.360 7.380 1.715 ;
        RECT  6.425 1.365 6.805 3.260 ;
        RECT  5.770 1.360 6.110 1.715 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.285 2.250 3.040 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.405 -0.400 6.745 1.135 ;
        RECT  5.170 -0.400 5.510 1.085 ;
        RECT  3.640 -0.400 3.980 1.040 ;
        RECT  1.685 -0.400 2.025 1.400 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.460 3.560 6.800 5.280 ;
        RECT  5.225 3.555 5.565 5.280 ;
        RECT  2.450 3.370 2.790 5.280 ;
        RECT  0.790 3.960 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.795 2.910 3.510 3.140 ;
        RECT  3.170 2.910 3.510 4.175 ;
        RECT  1.795 2.910 2.070 4.185 ;
        RECT  1.730 3.840 2.070 4.185 ;
        RECT  0.945 1.060 1.300 2.020 ;
        RECT  0.945 1.790 3.700 2.020 ;
        RECT  3.355 1.790 3.700 2.130 ;
        RECT  0.945 1.060 1.285 2.985 ;
        RECT  2.870 0.840 3.225 1.560 ;
        RECT  2.870 1.270 4.230 1.560 ;
        RECT  3.930 2.120 4.420 2.460 ;
        RECT  3.930 1.270 4.230 4.180 ;
        RECT  3.890 2.810 4.230 4.180 ;
        RECT  4.590 1.360 4.930 1.700 ;
        RECT  4.650 1.945 5.870 2.285 ;
        RECT  4.650 1.360 4.930 3.260 ;
        RECT  4.590 2.915 4.930 3.260 ;
        RECT  0.945 1.790 2.20 2.020 ;
    END
END EO2X4

MACRO EO2X2
    CLASS CORE ;
    FOREIGN EO2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.640 6.240 3.560 ;
        RECT  6.010 1.250 6.240 3.560 ;
        RECT  5.850 1.250 6.240 1.590 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.285 2.250 3.040 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.418  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 0.720 ;
        RECT  5.290 -0.400 5.630 0.720 ;
        RECT  3.930 -0.400 4.270 1.040 ;
        RECT  1.805 -0.400 2.145 1.400 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.960 6.750 5.280 ;
        RECT  5.290 3.960 5.630 5.280 ;
        RECT  2.450 3.555 2.790 5.280 ;
        RECT  0.790 3.960 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.795 2.910 3.510 3.140 ;
        RECT  3.170 2.910 3.510 4.025 ;
        RECT  1.795 2.910 2.070 4.185 ;
        RECT  1.730 3.840 2.070 4.185 ;
        RECT  0.945 1.060 1.300 2.020 ;
        RECT  0.945 1.790 3.700 2.020 ;
        RECT  3.355 1.790 3.700 2.130 ;
        RECT  0.945 1.060 1.285 2.985 ;
        RECT  3.120 1.060 3.475 1.560 ;
        RECT  3.120 1.270 4.230 1.560 ;
        RECT  3.930 1.945 4.420 2.285 ;
        RECT  3.930 1.270 4.230 4.180 ;
        RECT  3.890 3.840 4.230 4.180 ;
        RECT  4.530 1.360 4.915 1.700 ;
        RECT  4.650 1.945 5.780 2.285 ;
        RECT  4.650 1.360 4.915 3.450 ;
        RECT  4.530 2.640 4.915 3.450 ;
        RECT  0.945 1.790 2.80 2.020 ;
    END
END EO2X2

MACRO EO2X1
    CLASS CORE ;
    FOREIGN EO2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.285 2.250 3.040 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.103  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 2.800 4.285 4.175 ;
        RECT  3.930 1.270 4.285 4.175 ;
        RECT  2.870 1.270 4.285 1.560 ;
        RECT  2.870 0.840 3.225 1.560 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  2.450 3.370 2.790 5.280 ;
        RECT  0.790 3.960 1.130 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.640 -0.400 3.980 1.040 ;
        RECT  1.685 -0.400 2.025 1.400 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.730 2.910 3.510 3.140 ;
        RECT  3.170 2.910 3.510 4.180 ;
        RECT  1.730 2.910 2.070 4.185 ;
        RECT  0.945 1.060 1.300 2.020 ;
        RECT  0.945 1.790 3.700 2.020 ;
        RECT  3.355 1.790 3.700 2.130 ;
        RECT  0.945 1.060 1.285 2.985 ;
        RECT  0.945 1.790 2.60 2.020 ;
    END
END EO2X1

MACRO EO2X0
    CLASS CORE ;
    FOREIGN EO2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.604  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.410 2.850 3.025 3.190 ;
        RECT  2.645 1.170 3.025 3.190 ;
        RECT  2.250 1.170 3.025 1.510 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.415 2.045 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.243  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.245 0.585 2.740 ;
        RECT  0.120 2.245 0.525 2.780 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.620 3.895 1.960 5.280 ;
        RECT  0.180 3.835 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.780 -0.400 2.590 0.710 ;
        RECT  0.180 -0.400 0.520 1.290 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.970 0.630 1.320 1.305 ;
        RECT  0.970 1.075 1.875 1.305 ;
        RECT  1.645 2.160 2.415 2.500 ;
        RECT  0.675 2.955 1.875 3.185 ;
        RECT  1.645 1.075 1.875 3.185 ;
        RECT  0.180 3.010 0.830 3.240 ;
        RECT  0.180 3.010 0.520 3.295 ;
        RECT  0.955 3.435 2.730 3.665 ;
        RECT  2.390 3.435 2.730 3.910 ;
        RECT  0.900 3.460 1.240 4.165 ;
    END
END EO2X0

MACRO EN3X4
    CLASS CORE ;
    FOREIGN EN3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.559  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.975 3.470 5.545 4.250 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 2.675 3.000 ;
        RECT  1.940 2.250 2.675 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.922  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.660 2.920 11.160 3.260 ;
        RECT  9.550 1.360 11.160 1.710 ;
        RECT  10.820 1.350 11.160 1.710 ;
        RECT  10.205 1.360 10.585 3.260 ;
        RECT  9.550 1.335 9.890 1.710 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.185 -0.400 10.525 1.130 ;
        RECT  8.950 -0.400 9.290 1.080 ;
        RECT  6.230 -0.400 6.570 1.340 ;
        RECT  3.575 -0.400 3.960 1.040 ;
        RECT  1.665 -0.400 2.005 1.340 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.240 3.560 10.580 5.280 ;
        RECT  9.005 3.555 9.345 5.280 ;
        RECT  7.670 3.070 8.010 5.280 ;
        RECT  5.785 2.820 6.150 5.280 ;
        RECT  4.435 2.820 4.715 5.280 ;
        RECT  4.325 2.820 4.715 3.160 ;
        RECT  2.425 3.825 2.765 5.280 ;
        RECT  0.560 3.960 0.900 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.945 1.000 1.300 2.020 ;
        RECT  0.945 1.790 3.345 2.020 ;
        RECT  3.000 1.790 3.345 2.130 ;
        RECT  0.945 1.000 1.285 2.985 ;
        RECT  1.705 3.355 3.485 3.585 ;
        RECT  3.145 3.355 3.485 4.150 ;
        RECT  1.705 3.355 2.045 4.185 ;
        RECT  4.315 0.630 4.910 0.940 ;
        RECT  2.805 1.000 3.160 1.560 ;
        RECT  4.315 0.630 4.580 1.560 ;
        RECT  2.805 1.270 4.580 1.560 ;
        RECT  3.865 1.270 4.095 4.180 ;
        RECT  3.865 3.820 4.205 4.180 ;
        RECT  5.510 1.000 5.850 1.800 ;
        RECT  6.950 1.000 7.290 1.800 ;
        RECT  5.510 1.570 7.290 1.800 ;
        RECT  4.810 1.170 5.150 2.370 ;
        RECT  4.810 2.030 7.480 2.370 ;
        RECT  5.035 2.030 5.375 3.160 ;
        RECT  7.670 1.000 8.010 1.340 ;
        RECT  7.725 1.000 8.010 2.455 ;
        RECT  7.725 2.115 8.295 2.455 ;
        RECT  7.725 1.000 8.000 2.830 ;
        RECT  6.950 2.600 8.000 2.830 ;
        RECT  6.950 2.600 7.290 3.880 ;
        RECT  8.370 1.355 8.755 1.695 ;
        RECT  8.525 1.940 9.650 2.280 ;
        RECT  8.525 1.355 8.755 3.260 ;
        RECT  8.370 2.915 8.755 3.260 ;
        RECT  0.945 1.790 2.60 2.020 ;
        RECT  4.810 2.030 6.90 2.370 ;
    END
END EN3X4

MACRO EN3X2
    CLASS CORE ;
    FOREIGN EN3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.367  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.975 3.470 5.545 4.250 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 2.675 3.000 ;
        RECT  1.940 2.250 2.675 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.640 10.030 3.560 ;
        RECT  9.790 1.250 10.030 3.560 ;
        RECT  9.630 1.250 10.030 1.590 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 0.720 ;
        RECT  9.070 -0.400 9.410 0.720 ;
        RECT  6.230 -0.400 6.570 1.340 ;
        RECT  3.575 -0.400 3.960 1.040 ;
        RECT  1.665 -0.400 2.005 1.340 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 3.960 10.530 5.280 ;
        RECT  9.070 3.960 9.410 5.280 ;
        RECT  7.670 3.840 8.010 5.280 ;
        RECT  5.775 2.820 6.150 5.280 ;
        RECT  4.435 2.820 4.715 5.280 ;
        RECT  4.325 2.820 4.715 3.160 ;
        RECT  2.425 3.825 2.765 5.280 ;
        RECT  0.560 3.960 0.900 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.945 1.000 1.300 2.020 ;
        RECT  0.945 1.790 3.345 2.020 ;
        RECT  3.000 1.790 3.345 2.130 ;
        RECT  0.945 1.000 1.285 2.985 ;
        RECT  1.705 3.355 3.485 3.585 ;
        RECT  3.145 3.355 3.485 4.150 ;
        RECT  1.705 3.355 2.045 4.185 ;
        RECT  4.315 0.630 4.910 0.940 ;
        RECT  2.805 1.000 3.160 1.560 ;
        RECT  4.315 0.630 4.580 1.560 ;
        RECT  2.805 1.270 4.580 1.560 ;
        RECT  3.865 1.270 4.095 4.180 ;
        RECT  3.865 3.820 4.205 4.180 ;
        RECT  5.510 1.000 5.850 1.800 ;
        RECT  6.950 1.000 7.290 1.800 ;
        RECT  5.510 1.570 7.290 1.800 ;
        RECT  4.810 1.170 5.150 2.370 ;
        RECT  4.810 2.030 7.480 2.370 ;
        RECT  5.035 2.030 5.375 3.160 ;
        RECT  7.710 1.945 8.290 2.285 ;
        RECT  7.710 1.360 8.050 2.830 ;
        RECT  6.950 2.600 8.050 2.830 ;
        RECT  6.950 2.600 7.290 4.180 ;
        RECT  8.270 0.665 8.750 1.005 ;
        RECT  8.520 1.945 9.560 2.285 ;
        RECT  8.520 0.665 8.750 3.560 ;
        RECT  8.310 2.640 8.750 3.560 ;
        RECT  0.945 1.790 2.80 2.020 ;
        RECT  4.810 2.030 6.20 2.370 ;
    END
END EN3X2

MACRO EN3X1
    CLASS CORE ;
    FOREIGN EN3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.046  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 2.600 8.065 2.830 ;
        RECT  7.685 1.360 8.065 2.830 ;
        RECT  6.950 2.600 7.290 3.870 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.565  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.975 3.470 5.545 4.250 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.550 2.255 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.330 2.250 2.675 3.000 ;
        RECT  1.940 2.250 2.675 2.630 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.230 -0.400 6.570 1.340 ;
        RECT  3.575 -0.400 3.960 1.040 ;
        RECT  1.665 -0.400 2.005 1.340 ;
        RECT  0.180 -0.400 0.520 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.670 3.060 8.010 5.280 ;
        RECT  5.785 2.820 6.150 5.280 ;
        RECT  4.435 2.820 4.715 5.280 ;
        RECT  4.325 2.820 4.715 3.160 ;
        RECT  2.425 3.825 2.765 5.280 ;
        RECT  0.560 3.960 0.900 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.945 1.000 1.300 2.020 ;
        RECT  0.945 1.790 3.345 2.020 ;
        RECT  3.000 1.790 3.345 2.130 ;
        RECT  0.945 1.000 1.285 2.985 ;
        RECT  1.705 3.355 3.485 3.585 ;
        RECT  3.145 3.355 3.485 4.150 ;
        RECT  1.705 3.355 2.045 4.185 ;
        RECT  4.315 0.630 4.910 0.940 ;
        RECT  2.805 1.000 3.160 1.560 ;
        RECT  4.315 0.630 4.580 1.560 ;
        RECT  2.805 1.270 4.580 1.560 ;
        RECT  3.865 1.270 4.095 4.180 ;
        RECT  3.865 3.820 4.205 4.180 ;
        RECT  5.510 1.000 5.850 1.800 ;
        RECT  6.950 1.360 7.290 1.800 ;
        RECT  5.510 1.570 7.290 1.800 ;
        RECT  4.810 1.170 5.150 2.370 ;
        RECT  4.810 2.030 7.455 2.370 ;
        RECT  5.035 2.030 5.375 3.160 ;
        RECT  0.945 1.790 2.80 2.020 ;
        RECT  4.810 2.030 6.30 2.370 ;
    END
END EN3X1

MACRO EN3X0
    CLASS CORE ;
    FOREIGN EN3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.490  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.345 2.530 5.545 2.760 ;
        RECT  5.165 1.360 5.545 2.760 ;
        RECT  4.945 1.360 5.545 1.700 ;
        RECT  4.345 2.530 4.685 3.140 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.266  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 1.640 3.655 2.545 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.209  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.755 1.930 2.395 2.285 ;
        RECT  2.015 1.640 2.395 2.285 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.209  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.020 3.025 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 2.990 5.490 5.280 ;
        RECT  4.345 3.530 4.685 5.280 ;
        RECT  2.730 2.860 3.070 5.280 ;
        RECT  1.130 3.680 1.470 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.185 -0.400 4.525 0.670 ;
        RECT  2.620 -0.400 2.960 1.540 ;
        RECT  0.550 -0.400 1.360 0.740 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.200 0.890 1.540 ;
        RECT  0.180 1.200 0.520 4.095 ;
        RECT  0.180 3.755 0.735 4.095 ;
        RECT  1.820 0.630 2.170 1.305 ;
        RECT  1.295 1.075 2.170 1.305 ;
        RECT  0.750 1.770 1.525 2.110 ;
        RECT  1.295 1.075 1.525 2.990 ;
        RECT  1.295 2.650 1.825 2.990 ;
        RECT  0.780 2.640 1.065 3.450 ;
        RECT  0.780 3.220 2.270 3.450 ;
        RECT  1.930 3.220 2.270 3.795 ;
        RECT  4.145 1.400 4.485 2.300 ;
        RECT  4.145 1.960 4.935 2.300 ;
        RECT  3.885 2.070 4.935 2.300 ;
        RECT  3.885 2.070 4.115 3.870 ;
        RECT  3.530 3.530 4.115 3.870 ;
        RECT  3.370 0.700 3.720 1.130 ;
        RECT  4.945 0.640 5.285 1.130 ;
        RECT  3.370 0.900 5.285 1.130 ;
    END
END EN3X0

MACRO EN2X4
    CLASS CORE ;
    FOREIGN EN2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.565  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.490 3.850 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.922  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.880 2.920 7.380 3.260 ;
        RECT  5.770 1.365 7.380 1.715 ;
        RECT  7.040 1.355 7.380 1.715 ;
        RECT  6.425 1.365 6.805 3.260 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.565  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.525 0.550 2.255 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.460 3.560 6.800 5.280 ;
        RECT  5.225 3.560 5.565 5.280 ;
        RECT  3.890 2.760 4.230 5.280 ;
        RECT  2.005 2.810 2.370 5.280 ;
        RECT  0.155 2.720 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.405 -0.400 6.745 1.135 ;
        RECT  5.170 -0.400 5.510 1.085 ;
        RECT  2.450 -0.400 2.790 1.040 ;
        RECT  0.180 -0.400 0.520 0.960 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.730 0.875 2.070 1.500 ;
        RECT  3.170 1.060 3.510 1.500 ;
        RECT  1.730 1.270 3.510 1.500 ;
        RECT  1.010 0.640 1.350 2.070 ;
        RECT  0.900 1.730 3.700 2.070 ;
        RECT  0.900 1.725 1.240 3.060 ;
        RECT  3.890 1.060 4.230 1.400 ;
        RECT  3.930 1.060 4.230 2.530 ;
        RECT  3.930 2.115 4.485 2.530 ;
        RECT  3.170 2.300 4.485 2.530 ;
        RECT  3.170 2.300 3.510 3.500 ;
        RECT  4.590 1.360 4.945 1.700 ;
        RECT  4.715 1.995 5.870 2.335 ;
        RECT  4.715 1.360 4.945 3.260 ;
        RECT  4.590 2.915 4.945 3.260 ;
        RECT  0.900 1.730 2.70 2.070 ;
    END
END EN2X4

MACRO EN2X2
    CLASS CORE ;
    FOREIGN EN2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.364  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.490 3.850 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.750 6.190 3.560 ;
        RECT  5.960 1.250 6.190 3.560 ;
        RECT  5.850 1.250 6.190 1.590 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.364  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.525 0.550 2.255 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.405 3.960 6.750 5.280 ;
        RECT  5.290 3.960 5.630 5.280 ;
        RECT  3.830 2.760 4.170 5.280 ;
        RECT  1.945 2.810 2.310 5.280 ;
        RECT  0.155 2.720 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 0.720 ;
        RECT  5.290 -0.400 5.630 0.720 ;
        RECT  2.450 -0.400 2.790 1.040 ;
        RECT  0.180 -0.400 0.520 0.960 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.730 0.700 2.070 1.500 ;
        RECT  3.170 0.700 3.510 1.500 ;
        RECT  1.730 1.270 3.510 1.500 ;
        RECT  1.010 0.640 1.350 2.070 ;
        RECT  0.900 1.730 3.700 2.070 ;
        RECT  0.900 1.725 1.240 3.060 ;
        RECT  3.890 0.700 4.230 1.040 ;
        RECT  3.930 0.700 4.230 2.285 ;
        RECT  3.930 1.945 4.425 2.285 ;
        RECT  3.930 0.700 4.220 2.530 ;
        RECT  3.110 2.300 4.220 2.530 ;
        RECT  3.110 2.300 3.450 3.060 ;
        RECT  4.490 1.360 4.915 1.700 ;
        RECT  4.655 1.945 5.725 2.285 ;
        RECT  4.655 1.360 4.915 3.560 ;
        RECT  4.530 2.750 4.915 3.560 ;
        RECT  0.900 1.730 2.30 2.070 ;
    END
END EN2X2

MACRO EN2X1
    CLASS CORE ;
    FOREIGN EN2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.562  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.490 3.850 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.046  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.170 2.300 4.285 2.530 ;
        RECT  3.905 1.060 4.285 2.530 ;
        RECT  3.890 1.060 4.285 1.400 ;
        RECT  3.170 2.300 3.510 3.500 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.562  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.525 0.550 2.255 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.890 2.760 4.230 5.280 ;
        RECT  2.005 2.640 2.370 5.280 ;
        RECT  0.155 2.720 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  2.450 -0.400 2.790 1.040 ;
        RECT  0.180 -0.400 0.520 0.960 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.730 0.875 2.070 1.500 ;
        RECT  3.170 1.060 3.510 1.500 ;
        RECT  1.730 1.270 3.510 1.500 ;
        RECT  1.010 0.640 1.350 2.070 ;
        RECT  0.900 1.730 3.675 2.070 ;
        RECT  0.900 1.725 1.240 3.060 ;
        RECT  0.900 1.730 2.70 2.070 ;
    END
END EN2X1

MACRO EN2X0
    CLASS CORE ;
    FOREIGN EN2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.360 3.025 2.020 ;
        RECT  1.865 3.005 2.975 3.310 ;
        RECT  2.645 1.360 2.975 3.310 ;
        RECT  2.425 1.360 3.025 1.700 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.266  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.975 1.430 2.315 ;
        RECT  0.755 1.975 1.135 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.266  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.620 0.525 2.220 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.090 3.840 2.900 5.280 ;
        RECT  0.490 2.980 0.830 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.660 -0.400 2.000 0.670 ;
        RECT  0.180 -0.400 0.520 1.040 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.625 1.400 1.970 1.740 ;
        RECT  1.660 1.400 1.970 2.775 ;
        RECT  1.660 2.420 2.415 2.775 ;
        RECT  1.400 2.545 2.415 2.775 ;
        RECT  1.400 2.545 1.630 4.180 ;
        RECT  1.290 3.840 1.630 4.180 ;
        RECT  0.890 0.700 1.240 1.130 ;
        RECT  2.425 0.640 2.765 1.130 ;
        RECT  0.890 0.900 2.765 1.130 ;
    END
END EN2X0

MACRO DLY8X1
    CLASS CORE ;
    FOREIGN DLY8X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 2.850 12.475 3.770 ;
        RECT  12.200 1.245 12.475 3.770 ;
        RECT  12.080 1.245 12.475 1.590 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.505 2.735 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.880 -0.400 11.820 0.750 ;
        RECT  7.070 -0.400 7.410 1.000 ;
        RECT  5.430 -0.400 5.770 0.750 ;
        RECT  0.510 -0.400 1.790 0.750 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.320 3.575 11.660 5.280 ;
        RECT  6.400 3.880 6.740 5.280 ;
        RECT  0.880 3.790 1.220 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.220 1.015 1.560 ;
        RECT  0.735 2.360 2.490 2.700 ;
        RECT  0.735 1.220 1.015 3.560 ;
        RECT  0.180 3.330 1.015 3.560 ;
        RECT  0.180 3.330 0.520 4.210 ;
        RECT  2.830 2.610 6.060 2.950 ;
        RECT  2.830 1.970 3.170 3.195 ;
        RECT  2.590 2.915 2.870 4.130 ;
        RECT  2.530 3.790 2.870 4.130 ;
        RECT  3.910 1.890 4.250 2.230 ;
        RECT  3.910 1.950 6.570 2.230 ;
        RECT  6.290 2.450 8.340 2.790 ;
        RECT  6.290 1.950 6.570 3.540 ;
        RECT  3.400 3.260 6.570 3.540 ;
        RECT  3.400 3.260 3.630 4.210 ;
        RECT  3.230 3.890 3.630 4.210 ;
        RECT  8.510 1.880 8.955 2.220 ;
        RECT  8.675 2.495 11.100 2.835 ;
        RECT  8.675 1.880 8.955 3.515 ;
        RECT  8.520 3.175 8.955 3.515 ;
        RECT  9.570 1.530 9.910 2.230 ;
        RECT  9.570 1.950 11.970 2.230 ;
        RECT  11.330 1.950 11.970 2.290 ;
        RECT  11.330 1.950 11.610 3.345 ;
        RECT  9.230 3.065 11.610 3.345 ;
        RECT  9.230 3.065 9.570 4.170 ;
        RECT  2.830 2.610 5.90 2.950 ;
        RECT  3.910 1.950 5.70 2.230 ;
        RECT  6.290 2.450 7.80 2.790 ;
        RECT  3.400 3.260 5.30 3.540 ;
        RECT  8.675 2.495 10.20 2.835 ;
        RECT  9.570 1.950 10.80 2.230 ;
        RECT  9.230 3.065 10.60 3.345 ;
    END
END DLY8X1

MACRO DLY8X0
    CLASS CORE ;
    FOREIGN DLY8X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 2.860 12.475 3.600 ;
        RECT  12.200 1.360 12.475 3.600 ;
        RECT  12.080 1.360 12.475 1.705 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.505 2.735 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.280 -0.400 11.620 1.700 ;
        RECT  10.680 -0.400 11.620 1.150 ;
        RECT  6.700 -0.400 7.040 1.000 ;
        RECT  5.430 -0.400 5.770 0.750 ;
        RECT  0.510 -0.400 1.790 0.750 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.480 3.910 11.820 5.280 ;
        RECT  6.380 3.160 6.720 5.280 ;
        RECT  0.880 3.790 1.220 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.110 1.015 1.450 ;
        RECT  0.735 2.360 2.490 2.700 ;
        RECT  0.735 1.110 1.015 3.560 ;
        RECT  0.180 3.330 1.015 3.560 ;
        RECT  0.180 3.330 0.520 4.110 ;
        RECT  2.830 1.970 3.170 2.950 ;
        RECT  2.830 2.610 5.630 2.950 ;
        RECT  2.830 1.970 3.110 4.095 ;
        RECT  2.710 3.755 3.110 4.095 ;
        RECT  7.430 0.660 8.370 1.000 ;
        RECT  3.910 1.890 4.250 2.230 ;
        RECT  3.910 1.950 6.140 2.230 ;
        RECT  5.860 2.450 8.460 2.790 ;
        RECT  5.860 1.950 6.140 4.170 ;
        RECT  3.410 3.890 6.140 4.170 ;
        RECT  3.410 3.890 3.750 4.230 ;
        RECT  9.380 0.910 10.320 1.250 ;
        RECT  8.140 1.880 8.970 2.220 ;
        RECT  8.690 2.610 11.100 2.950 ;
        RECT  8.690 1.880 8.970 4.180 ;
        RECT  8.500 3.840 8.970 4.180 ;
        RECT  9.370 1.880 9.710 2.230 ;
        RECT  9.370 1.950 11.970 2.230 ;
        RECT  11.330 1.950 11.970 2.290 ;
        RECT  11.330 1.950 11.610 3.540 ;
        RECT  9.200 3.260 11.610 3.540 ;
        RECT  9.200 3.260 9.540 4.080 ;
        RECT  2.830 2.610 4.40 2.950 ;
        RECT  3.910 1.950 5.90 2.230 ;
        RECT  5.860 2.450 7.40 2.790 ;
        RECT  3.410 3.890 5.60 4.170 ;
        RECT  8.690 2.610 10.50 2.950 ;
        RECT  9.370 1.950 10.30 2.230 ;
        RECT  9.200 3.260 10.40 3.540 ;
    END
END DLY8X0

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.000 2.860 7.435 3.885 ;
        RECT  7.155 1.245 7.435 3.885 ;
        RECT  7.000 1.245 7.435 1.590 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.505 2.735 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.240 -0.400 6.580 1.700 ;
        RECT  5.430 -0.400 6.580 0.750 ;
        RECT  0.980 -0.400 1.790 0.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.230 3.770 6.570 5.280 ;
        RECT  0.880 3.790 1.220 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.220 1.015 1.560 ;
        RECT  0.735 2.360 2.490 2.700 ;
        RECT  0.735 1.220 1.015 3.560 ;
        RECT  0.180 3.330 1.015 3.560 ;
        RECT  0.180 3.330 0.520 4.210 ;
        RECT  2.830 2.610 6.060 2.950 ;
        RECT  2.830 1.970 3.170 3.590 ;
        RECT  2.730 3.250 3.170 3.590 ;
        RECT  3.910 1.690 4.250 2.230 ;
        RECT  3.910 1.950 6.860 2.230 ;
        RECT  6.290 1.950 6.860 2.290 ;
        RECT  6.290 1.950 6.570 3.540 ;
        RECT  3.520 3.260 6.570 3.540 ;
        RECT  3.520 3.260 3.860 3.600 ;
        RECT  2.830 2.610 5.60 2.950 ;
        RECT  3.910 1.950 5.50 2.230 ;
        RECT  3.520 3.260 5.20 3.540 ;
    END
END DLY4X1

MACRO DLY4X0
    CLASS CORE ;
    FOREIGN DLY4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.637  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 3.910 7.435 4.250 ;
        RECT  7.155 1.360 7.435 4.250 ;
        RECT  7.055 2.860 7.435 3.240 ;
        RECT  7.040 1.360 7.435 1.705 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.505 2.735 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.240 -0.400 6.580 1.700 ;
        RECT  5.430 -0.400 6.580 0.955 ;
        RECT  0.510 -0.400 1.790 0.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 3.930 6.660 5.280 ;
        RECT  0.880 3.790 1.220 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.250 1.015 1.590 ;
        RECT  0.735 2.360 2.490 2.700 ;
        RECT  0.735 1.250 1.015 3.560 ;
        RECT  0.180 3.330 1.015 3.560 ;
        RECT  0.180 3.330 0.520 4.115 ;
        RECT  3.920 0.655 5.060 0.995 ;
        RECT  2.830 2.610 6.060 2.950 ;
        RECT  2.830 1.970 3.170 3.195 ;
        RECT  2.590 2.915 2.870 4.130 ;
        RECT  2.530 3.790 2.870 4.130 ;
        RECT  3.910 1.890 4.250 2.230 ;
        RECT  3.910 1.950 6.925 2.230 ;
        RECT  2.830 2.610 5.60 2.950 ;
        RECT  3.910 1.950 5.40 2.230 ;
        RECT  6.290 1.950 6.925 2.290 ;
        RECT  6.290 1.950 6.570 3.700 ;
        RECT  3.320 3.420 6.570 3.700 ;
        RECT  3.320 3.420 3.660 3.760 ;
    END
END DLY4X0

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.740 2.860 6.175 3.885 ;
        RECT  5.895 1.245 6.175 3.885 ;
        RECT  5.740 1.245 6.175 1.590 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.505 2.735 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.980 -0.400 5.320 1.700 ;
        RECT  0.780 -0.400 1.120 0.750 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.970 3.770 5.310 5.280 ;
        RECT  0.940 3.790 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.220 1.015 1.560 ;
        RECT  0.735 2.545 2.070 2.885 ;
        RECT  0.735 1.220 1.015 3.425 ;
        RECT  0.180 3.085 1.015 3.425 ;
        RECT  2.235 1.970 2.540 2.310 ;
        RECT  2.300 1.970 2.540 3.590 ;
        RECT  2.300 2.610 4.715 2.950 ;
        RECT  2.300 2.610 2.570 3.590 ;
        RECT  2.230 3.255 2.570 3.590 ;
        RECT  3.420 1.690 3.760 2.230 ;
        RECT  3.420 1.950 5.600 2.230 ;
        RECT  5.045 1.950 5.600 2.395 ;
        RECT  5.045 1.950 5.325 3.540 ;
        RECT  3.125 3.260 5.325 3.540 ;
        RECT  3.125 3.260 3.465 3.600 ;
        RECT  2.300 2.610 3.80 2.950 ;
        RECT  3.420 1.950 4.80 2.230 ;
        RECT  3.125 3.260 4.70 3.540 ;
    END
END DLY2X1

MACRO DLY2X0
    CLASS CORE ;
    FOREIGN DLY2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.040 2.740 5.545 3.240 ;
        RECT  5.265 1.330 5.545 3.240 ;
        RECT  5.150 1.330 5.545 1.675 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.530 0.505 3.240 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.145 -0.400 5.485 0.875 ;
        RECT  4.280 -0.400 4.625 1.050 ;
        RECT  0.905 -0.400 1.245 1.700 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.035 3.540 5.375 5.280 ;
        RECT  4.235 3.840 4.575 5.280 ;
        RECT  1.025 3.930 1.365 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.755 0.520 1.155 ;
        RECT  0.240 0.755 0.520 2.300 ;
        RECT  0.240 2.020 1.015 2.300 ;
        RECT  0.735 2.465 2.165 2.805 ;
        RECT  0.735 2.020 1.015 3.700 ;
        RECT  0.180 3.470 1.015 3.700 ;
        RECT  0.180 3.470 0.520 3.810 ;
        RECT  3.015 3.250 3.355 4.180 ;
        RECT  3.105 0.710 3.445 1.750 ;
        RECT  2.395 1.970 2.735 2.310 ;
        RECT  2.415 2.100 4.055 2.380 ;
        RECT  3.715 2.100 4.055 2.910 ;
        RECT  2.415 1.970 2.685 3.590 ;
        RECT  2.315 3.250 2.685 3.590 ;
        RECT  4.325 1.410 4.640 2.400 ;
        RECT  4.325 2.060 4.925 2.400 ;
        RECT  4.325 1.410 4.625 3.480 ;
        RECT  4.195 3.140 4.625 3.480 ;
    END
END DLY2X0

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.149  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.750 3.890 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.823  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 1.175 4.915 2.640 ;
        RECT  4.440 2.870 4.785 3.795 ;
        RECT  4.520 1.175 4.785 3.795 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.715 -0.400 4.060 1.265 ;
        RECT  0.980 -0.400 1.320 1.620 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.720 2.985 4.060 5.280 ;
        RECT  0.980 2.840 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.280 0.520 2.610 ;
        RECT  1.485 1.800 1.825 2.610 ;
        RECT  0.180 2.380 1.825 2.610 ;
        RECT  0.220 2.380 0.560 3.165 ;
        RECT  2.085 0.700 2.425 2.295 ;
        RECT  2.085 1.955 3.540 2.295 ;
        RECT  2.085 0.700 2.315 3.160 ;
        RECT  1.970 2.820 2.315 3.160 ;
        RECT  2.800 0.740 3.140 1.080 ;
        RECT  2.910 0.740 3.140 1.725 ;
        RECT  2.910 1.495 4.110 1.725 ;
        RECT  3.770 2.000 4.290 2.340 ;
        RECT  3.770 1.495 4.110 2.755 ;
        RECT  2.820 2.525 4.110 2.755 ;
        RECT  2.820 2.525 3.160 3.215 ;
    END
END DLY1X1

MACRO DLY1X0
    CLASS CORE ;
    FOREIGN DLY1X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.750 3.890 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 1.280 4.915 3.130 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.715 -0.400 4.060 1.265 ;
        RECT  0.810 -0.400 1.150 1.010 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.720 2.985 4.060 5.280 ;
        RECT  0.980 2.840 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.455 1.800 1.795 2.610 ;
        RECT  0.180 2.380 1.795 2.610 ;
        RECT  0.180 1.280 0.520 3.130 ;
        RECT  2.060 1.955 3.500 2.295 ;
        RECT  2.060 0.700 2.400 3.160 ;
        RECT  2.800 0.630 3.140 0.970 ;
        RECT  2.910 0.630 3.140 1.725 ;
        RECT  2.910 1.495 4.290 1.725 ;
        RECT  3.950 1.495 4.290 2.755 ;
        RECT  2.950 2.525 4.290 2.755 ;
        RECT  2.950 2.525 3.180 3.670 ;
        RECT  2.840 3.330 3.180 3.670 ;
    END
END DLY1X0

MACRO DLLX4
    CLASS CORE ;
    FOREIGN DLLX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.820 1.240 11.215 4.100 ;
        RECT  9.660 2.250 11.215 2.480 ;
        RECT  9.500 2.640 9.890 3.770 ;
        RECT  9.660 0.790 9.890 3.770 ;
        RECT  9.500 0.790 9.890 1.700 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.550 1.135 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.180 1.240 8.520 3.450 ;
        RECT  6.860 2.250 8.520 2.630 ;
        RECT  6.860 1.240 7.200 3.450 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.260 -0.400 10.600 0.720 ;
        RECT  6.100 -0.400 9.080 0.720 ;
        RECT  4.780 -0.400 5.120 0.985 ;
        RECT  2.460 -0.400 2.800 0.955 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  6.300 4.140 10.400 5.280 ;
        RECT  4.780 4.150 5.120 5.280 ;
        RECT  2.205 3.785 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  1.330 2.145 1.670 2.480 ;
        RECT  1.340 2.125 1.670 2.480 ;
        RECT  0.180 2.250 1.670 2.480 ;
        RECT  0.180 2.250 0.520 3.460 ;
        RECT  3.875 2.455 4.215 3.460 ;
        RECT  0.180 3.230 4.215 3.460 ;
        RECT  1.700 0.980 2.130 1.320 ;
        RECT  3.940 1.785 4.225 2.125 ;
        RECT  3.315 1.895 4.225 2.125 ;
        RECT  1.740 2.700 2.130 3.000 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.710 2.130 3.000 ;
        RECT  3.155 2.700 3.545 3.000 ;
        RECT  3.315 1.895 3.545 3.000 ;
        RECT  1.700 2.770 3.545 3.000 ;
        RECT  3.660 1.215 4.000 1.555 ;
        RECT  3.660 1.325 4.685 1.555 ;
        RECT  4.455 1.880 6.120 2.110 ;
        RECT  5.780 1.880 6.120 2.220 ;
        RECT  4.455 1.325 4.685 3.920 ;
        RECT  3.435 3.690 4.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  5.540 1.240 6.630 1.580 ;
        RECT  8.895 2.075 9.430 2.415 ;
        RECT  4.915 2.340 5.235 2.680 ;
        RECT  4.915 2.450 6.630 2.680 ;
        RECT  6.400 1.240 6.630 3.910 ;
        RECT  8.895 2.075 9.125 3.910 ;
        RECT  6.400 3.680 9.125 3.910 ;
        RECT  5.540 2.450 5.880 4.170 ;
        RECT  0.180 3.230 3.00 3.460 ;
        RECT  6.400 3.680 8.60 3.910 ;
    END
END DLLX4

MACRO DLLX2
    CLASS CORE ;
    FOREIGN DLLX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.240 1.135 3.480 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.785 1.615 6.445 2.080 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.550 8.175 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.240 2.400 3.480 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.320 ;
        RECT  6.160 -0.400 6.500 0.850 ;
        RECT  4.190 -0.400 4.530 0.810 ;
        RECT  2.820 -0.400 3.160 0.720 ;
        RECT  0.180 -0.400 1.640 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.740 3.950 8.080 5.280 ;
        RECT  6.370 3.750 6.710 5.280 ;
        RECT  3.700 3.910 4.045 5.280 ;
        RECT  1.500 4.170 2.960 5.280 ;
        RECT  0.180 4.010 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.190 1.240 3.720 1.580 ;
        RECT  3.190 2.690 4.045 3.030 ;
        RECT  3.190 2.690 3.720 3.550 ;
        RECT  3.190 1.240 3.420 3.940 ;
        RECT  0.930 3.710 3.420 3.940 ;
        RECT  0.930 3.710 1.270 4.070 ;
        RECT  5.130 0.630 5.470 1.415 ;
        RECT  4.275 1.180 5.470 1.415 ;
        RECT  3.650 2.020 4.505 2.360 ;
        RECT  4.275 1.180 4.505 4.035 ;
        RECT  4.275 3.750 5.480 4.035 ;
        RECT  6.690 0.990 7.200 1.330 ;
        RECT  4.850 1.680 5.555 2.020 ;
        RECT  5.325 1.680 5.555 3.060 ;
        RECT  6.690 0.990 6.920 3.060 ;
        RECT  5.325 2.720 5.760 3.060 ;
        RECT  6.690 2.720 7.250 3.060 ;
        RECT  5.325 2.830 7.250 3.060 ;
        RECT  8.300 0.980 8.640 1.320 ;
        RECT  7.150 2.125 7.480 2.480 ;
        RECT  7.150 2.145 7.490 2.480 ;
        RECT  7.150 2.250 8.640 2.480 ;
        RECT  4.750 2.350 5.090 3.520 ;
        RECT  8.300 2.250 8.640 3.520 ;
        RECT  8.405 0.980 8.640 3.520 ;
        RECT  4.750 3.290 8.640 3.520 ;
        RECT  0.930 3.710 2.50 3.940 ;
        RECT  4.750 3.290 7.60 3.520 ;
    END
END DLLX2

MACRO DLLX1
    CLASS CORE ;
    FOREIGN DLLX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.820 0.520 3.880 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 2.970 1.960 3.780 ;
        RECT  1.620 0.700 1.960 1.040 ;
        RECT  1.620 0.700 1.850 1.495 ;
        RECT  1.385 2.250 1.765 2.630 ;
        RECT  1.470 1.265 1.700 3.215 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.840 2.095 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.500 7.530 1.840 ;
        RECT  7.055 1.500 7.435 2.635 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.945 -0.400 7.285 1.270 ;
        RECT  5.525 -0.400 5.865 1.375 ;
        RECT  2.425 -0.400 3.235 0.710 ;
        RECT  0.900 -0.400 1.240 1.060 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.910 3.525 7.250 5.280 ;
        RECT  5.810 3.800 6.150 5.280 ;
        RECT  3.095 3.530 3.500 5.280 ;
        RECT  0.900 3.030 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.160 1.360 2.500 1.700 ;
        RECT  2.160 1.360 2.425 2.350 ;
        RECT  1.995 2.010 2.425 2.350 ;
        RECT  2.195 1.360 2.425 3.850 ;
        RECT  2.195 3.510 2.715 3.850 ;
        RECT  3.440 1.035 4.465 1.375 ;
        RECT  3.440 1.035 3.670 2.780 ;
        RECT  2.655 2.440 3.670 2.780 ;
        RECT  2.655 2.480 3.960 2.780 ;
        RECT  3.730 2.480 3.960 3.940 ;
        RECT  3.730 3.600 4.790 3.940 ;
        RECT  6.110 0.810 6.565 1.155 ;
        RECT  3.900 1.605 4.915 1.945 ;
        RECT  4.685 1.605 4.915 2.835 ;
        RECT  4.685 2.415 5.200 2.835 ;
        RECT  6.110 0.810 6.340 2.835 ;
        RECT  4.685 2.550 6.340 2.835 ;
        RECT  7.665 0.865 8.010 1.205 ;
        RECT  6.570 1.980 6.825 3.295 ;
        RECT  7.660 2.820 8.010 3.295 ;
        RECT  7.775 0.865 8.010 3.295 ;
        RECT  4.190 3.065 8.010 3.295 ;
        RECT  4.190 3.010 4.530 3.350 ;
        RECT  4.190 3.065 7.60 3.295 ;
    END
END DLLX1

MACRO DLLX0
    CLASS CORE ;
    FOREIGN DLLX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.559  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.130 0.815 3.470 ;
        RECT  0.125 0.630 0.520 3.470 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.545  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.885 1.640 2.395 2.020 ;
        RECT  1.775 2.840 2.115 3.180 ;
        RECT  1.885 1.415 2.115 3.180 ;
        RECT  1.680 1.415 2.115 1.700 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.345 3.240 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.230 6.245 2.755 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.310 -0.400 6.650 1.090 ;
        RECT  4.910 -0.400 5.250 1.590 ;
        RECT  2.480 -0.400 2.820 0.970 ;
        RECT  0.880 -0.400 1.220 0.725 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.520 3.965 6.590 5.280 ;
        RECT  2.805 3.470 3.145 5.280 ;
        RECT  0.475 3.930 0.815 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.680 0.630 2.020 1.185 ;
        RECT  1.220 0.955 2.020 1.185 ;
        RECT  1.220 0.955 1.450 2.510 ;
        RECT  1.050 2.170 1.655 2.510 ;
        RECT  1.050 2.170 1.280 4.250 ;
        RECT  1.050 3.980 1.615 4.250 ;
        RECT  2.770 1.200 3.850 1.540 ;
        RECT  2.770 1.200 3.000 3.240 ;
        RECT  2.345 3.010 3.770 3.240 ;
        RECT  2.345 3.010 2.575 3.750 ;
        RECT  1.510 3.410 2.575 3.750 ;
        RECT  3.540 3.010 3.770 4.250 ;
        RECT  3.540 3.965 4.280 4.250 ;
        RECT  5.610 0.630 5.950 2.000 ;
        RECT  5.610 1.770 6.865 2.000 ;
        RECT  6.560 1.770 6.865 2.365 ;
        RECT  6.560 1.770 6.790 3.275 ;
        RECT  5.650 2.985 6.790 3.275 ;
        RECT  7.070 1.360 7.380 1.665 ;
        RECT  3.230 1.770 3.570 2.540 ;
        RECT  3.230 2.200 4.800 2.540 ;
        RECT  4.075 2.200 4.305 3.735 ;
        RECT  7.040 3.140 7.380 3.735 ;
        RECT  7.095 1.360 7.380 3.735 ;
        RECT  4.075 3.505 7.380 3.735 ;
        RECT  4.075 3.505 6.30 3.735 ;
    END
END DLLX0

MACRO DLLSX4
    CLASS CORE ;
    FOREIGN DLLSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.580 1.610 6.175 2.020 ;
        END
    END GN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.070 1.240 10.410 3.450 ;
        RECT  8.750 2.250 10.410 2.630 ;
        RECT  8.750 1.240 9.090 3.450 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.805 1.640 4.285 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 1.240 13.105 4.100 ;
        RECT  11.550 2.250 13.105 2.480 ;
        RECT  11.390 2.640 11.780 3.770 ;
        RECT  11.550 0.790 11.780 3.770 ;
        RECT  11.390 0.790 11.780 1.700 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  12.150 -0.400 12.490 0.720 ;
        RECT  9.510 -0.400 10.970 0.720 ;
        RECT  6.870 -0.400 8.330 0.720 ;
        RECT  5.450 -0.400 5.790 1.380 ;
        RECT  4.030 -0.400 4.370 0.970 ;
        RECT  1.770 -0.400 2.110 0.950 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  10.830 4.170 12.290 5.280 ;
        RECT  7.990 4.140 9.850 5.280 ;
        RECT  6.710 2.705 7.050 5.280 ;
        RECT  5.170 3.625 5.510 5.280 ;
        RECT  3.925 3.900 4.265 5.280 ;
        RECT  1.540 4.110 1.880 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.875 1.410 ;
        RECT  1.535 1.180 1.875 2.090 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  2.110 1.235 3.140 1.575 ;
        RECT  2.110 1.235 2.340 2.550 ;
        RECT  1.845 2.320 2.340 2.550 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.845 2.320 2.075 3.610 ;
        RECT  0.170 3.380 2.340 3.610 ;
        RECT  2.110 3.380 2.340 3.855 ;
        RECT  2.110 3.625 3.035 3.855 ;
        RECT  2.695 3.625 3.035 3.965 ;
        RECT  4.730 1.040 5.070 1.380 ;
        RECT  4.520 1.150 4.750 2.935 ;
        RECT  3.030 2.595 4.750 2.935 ;
        RECT  6.170 1.040 6.640 1.380 ;
        RECT  3.235 1.805 3.575 2.145 ;
        RECT  2.570 1.915 3.575 2.145 ;
        RECT  4.980 2.080 5.310 2.480 ;
        RECT  6.405 1.040 6.640 2.480 ;
        RECT  4.980 2.250 6.640 2.480 ;
        RECT  2.305 2.780 2.800 3.080 ;
        RECT  2.570 1.915 2.800 3.395 ;
        RECT  2.570 3.165 6.270 3.395 ;
        RECT  5.930 2.250 6.270 3.550 ;
        RECT  10.785 2.075 11.320 2.415 ;
        RECT  7.430 1.240 7.770 3.910 ;
        RECT  10.785 2.075 11.015 3.910 ;
        RECT  7.430 3.680 11.015 3.910 ;
        RECT  0.170 3.380 1.20 3.610 ;
        RECT  2.570 3.165 5.40 3.395 ;
        RECT  7.430 3.680 10.80 3.910 ;
    END
END DLLSX4

MACRO DLLSX2
    CLASS CORE ;
    FOREIGN DLLSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 1.240 8.065 3.480 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.795 2.130 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 1.640 1.135 2.465 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 1.240 9.340 3.480 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.075 1.585 5.645 2.020 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  6.920 -0.400 9.900 0.720 ;
        RECT  4.940 -0.400 5.280 1.320 ;
        RECT  3.445 -0.400 3.785 0.955 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.560 4.010 9.900 5.280 ;
        RECT  7.120 4.170 8.580 5.280 ;
        RECT  5.025 3.700 5.365 5.280 ;
        RECT  3.850 3.875 4.190 5.280 ;
        RECT  1.440 4.170 1.780 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.950 ;
        RECT  0.180 0.630 0.410 2.925 ;
        RECT  1.365 1.890 1.650 2.925 ;
        RECT  0.180 2.695 1.650 2.925 ;
        RECT  0.740 2.695 1.080 3.150 ;
        RECT  1.880 1.270 2.585 1.610 ;
        RECT  0.170 3.155 0.510 3.610 ;
        RECT  0.170 3.380 2.110 3.610 ;
        RECT  1.880 1.270 2.110 3.935 ;
        RECT  1.880 3.705 2.960 3.935 ;
        RECT  2.620 3.705 2.960 4.240 ;
        RECT  1.965 0.680 3.045 1.020 ;
        RECT  4.025 0.980 4.560 1.320 ;
        RECT  2.815 0.680 3.045 3.010 ;
        RECT  4.025 0.980 4.255 3.010 ;
        RECT  2.815 2.670 3.240 3.010 ;
        RECT  4.025 2.710 4.605 3.010 ;
        RECT  2.815 2.780 4.605 3.010 ;
        RECT  5.660 0.980 6.125 1.320 ;
        RECT  4.505 2.080 4.845 2.480 ;
        RECT  4.505 2.250 6.125 2.480 ;
        RECT  2.340 2.090 2.585 3.470 ;
        RECT  5.785 2.250 6.125 3.470 ;
        RECT  5.890 0.980 6.125 3.470 ;
        RECT  2.340 3.240 6.125 3.470 ;
        RECT  6.360 1.170 6.700 3.940 ;
        RECT  6.360 3.710 9.150 3.940 ;
        RECT  8.810 3.710 9.150 4.070 ;
        RECT  2.340 3.240 5.40 3.470 ;
        RECT  6.360 3.710 8.90 3.940 ;
    END
END DLLSX2

MACRO DLLSX1
    CLASS CORE ;
    FOREIGN DLLSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.235 2.250 8.695 2.630 ;
        RECT  8.120 3.270 8.465 4.080 ;
        RECT  8.235 0.700 8.465 4.080 ;
        RECT  8.120 0.700 8.465 1.040 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.560 0.820 9.955 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.655 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.860 2.030 3.260 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.035 1.500 6.375 1.840 ;
        RECT  6.035 1.020 6.325 1.840 ;
        RECT  5.795 1.020 6.325 1.415 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.840 -0.400 9.180 1.060 ;
        RECT  7.320 -0.400 7.660 0.710 ;
        RECT  5.665 -0.400 6.005 0.710 ;
        RECT  4.165 -0.400 4.505 1.410 ;
        RECT  1.480 -0.400 1.820 1.180 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.840 3.330 9.180 5.280 ;
        RECT  7.185 4.170 7.525 5.280 ;
        RECT  5.885 3.525 6.225 5.280 ;
        RECT  4.570 3.525 4.910 5.280 ;
        RECT  1.750 3.840 2.095 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 1.210 0.520 1.640 ;
        RECT  0.170 1.410 2.155 1.640 ;
        RECT  1.815 1.410 2.155 1.895 ;
        RECT  0.170 1.210 0.400 3.250 ;
        RECT  0.170 3.020 1.120 3.250 ;
        RECT  0.890 3.020 1.120 4.175 ;
        RECT  0.890 3.835 1.280 4.175 ;
        RECT  2.430 1.250 3.105 1.590 ;
        RECT  0.630 2.155 0.970 2.495 ;
        RECT  0.630 2.230 2.660 2.495 ;
        RECT  2.430 1.250 2.660 3.755 ;
        RECT  2.430 3.525 3.510 3.755 ;
        RECT  3.170 3.525 3.510 3.845 ;
        RECT  2.485 0.630 3.675 0.970 ;
        RECT  4.885 0.810 5.245 1.150 ;
        RECT  3.445 0.630 3.675 2.835 ;
        RECT  4.885 0.810 5.115 2.835 ;
        RECT  3.445 2.470 3.920 2.835 ;
        RECT  4.885 2.550 5.410 2.835 ;
        RECT  3.445 2.605 5.410 2.835 ;
        RECT  6.600 0.980 6.985 1.320 ;
        RECT  5.345 1.760 5.630 2.320 ;
        RECT  5.345 2.075 6.985 2.320 ;
        RECT  2.890 2.680 3.215 3.295 ;
        RECT  6.635 0.980 6.985 3.295 ;
        RECT  2.890 3.065 6.985 3.295 ;
        RECT  7.300 1.170 7.750 1.510 ;
        RECT  7.300 2.130 7.985 2.505 ;
        RECT  7.300 1.170 7.530 3.820 ;
        RECT  7.185 3.445 7.530 3.820 ;
        RECT  0.630 2.230 1.50 2.495 ;
        RECT  2.890 3.065 5.60 3.295 ;
    END
END DLLSX1

MACRO DLLSX0
    CLASS CORE ;
    FOREIGN DLLSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.595 2.250 7.435 2.630 ;
        RECT  6.595 0.675 7.240 1.015 ;
        RECT  6.180 3.965 6.825 4.250 ;
        RECT  6.595 0.675 6.825 4.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.559  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 0.630 8.705 4.135 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.460 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.760 1.765 3.350 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.930 2.230 5.270 2.755 ;
        RECT  4.535 2.230 5.270 2.630 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.595 -0.400 7.940 0.970 ;
        RECT  5.450 -0.400 6.365 1.145 ;
        RECT  3.950 -0.400 4.290 1.540 ;
        RECT  1.320 -0.400 1.660 1.460 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.055 3.885 7.865 5.280 ;
        RECT  4.560 3.965 5.630 5.280 ;
        RECT  1.755 3.580 2.095 5.280 ;
        RECT  0.180 3.930 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.960 ;
        RECT  0.115 1.730 1.765 1.960 ;
        RECT  1.480 1.730 1.765 2.070 ;
        RECT  0.115 0.630 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  1.995 1.230 2.890 1.540 ;
        RECT  0.575 2.300 2.225 2.530 ;
        RECT  0.575 2.300 0.915 2.955 ;
        RECT  1.995 1.230 2.225 3.240 ;
        RECT  1.995 3.010 2.810 3.240 ;
        RECT  2.580 3.010 2.810 4.250 ;
        RECT  2.580 3.930 3.320 4.250 ;
        RECT  4.560 0.780 4.990 1.120 ;
        RECT  4.650 0.780 4.990 1.725 ;
        RECT  4.650 1.495 5.905 1.725 ;
        RECT  5.600 1.495 5.905 2.365 ;
        RECT  5.600 1.495 5.830 3.275 ;
        RECT  4.690 2.985 5.830 3.275 ;
        RECT  2.455 1.770 2.740 2.580 ;
        RECT  2.455 2.350 3.840 2.580 ;
        RECT  3.445 2.350 3.840 2.635 ;
        RECT  3.445 2.350 3.800 2.655 ;
        RECT  3.445 2.350 3.675 3.735 ;
        RECT  6.080 3.140 6.365 3.735 ;
        RECT  6.135 1.505 6.365 3.735 ;
        RECT  3.445 3.505 6.365 3.735 ;
        RECT  7.055 1.375 7.895 1.715 ;
        RECT  7.665 2.395 8.005 2.735 ;
        RECT  7.665 1.375 7.895 3.335 ;
        RECT  7.125 2.995 7.895 3.335 ;
        RECT  3.445 3.505 5.80 3.735 ;
    END
END DLLSX0

MACRO DLLSQX4
    CLASS CORE ;
    FOREIGN DLLSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.580 1.610 6.175 2.020 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.805 1.640 4.285 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 1.130 10.585 3.880 ;
        RECT  8.910 2.130 10.585 2.360 ;
        RECT  8.750 2.640 9.140 3.880 ;
        RECT  8.910 1.130 9.140 3.880 ;
        RECT  8.750 1.130 9.140 1.470 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.470 ;
        RECT  6.870 -0.400 8.330 0.720 ;
        RECT  5.450 -0.400 5.790 1.380 ;
        RECT  4.030 -0.400 4.370 0.970 ;
        RECT  1.770 -0.400 2.110 0.950 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 2.640 9.810 5.280 ;
        RECT  7.990 3.950 8.330 5.280 ;
        RECT  6.710 2.700 7.050 5.280 ;
        RECT  5.170 3.625 5.510 5.280 ;
        RECT  3.925 3.900 4.265 5.280 ;
        RECT  1.540 4.110 1.880 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.875 1.410 ;
        RECT  1.535 1.180 1.875 2.090 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  2.110 1.235 3.140 1.575 ;
        RECT  2.110 1.235 2.340 2.550 ;
        RECT  1.845 2.320 2.340 2.550 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.845 2.320 2.075 3.610 ;
        RECT  0.170 3.380 2.340 3.610 ;
        RECT  2.110 3.380 2.340 3.855 ;
        RECT  2.110 3.625 3.035 3.855 ;
        RECT  2.695 3.625 3.035 3.965 ;
        RECT  4.730 1.040 5.070 1.380 ;
        RECT  4.520 1.150 4.750 2.935 ;
        RECT  3.030 2.595 4.750 2.935 ;
        RECT  6.170 1.040 6.640 1.380 ;
        RECT  3.235 1.805 3.575 2.145 ;
        RECT  2.570 1.915 3.575 2.145 ;
        RECT  4.980 2.080 5.310 2.480 ;
        RECT  6.405 1.040 6.640 2.480 ;
        RECT  4.980 2.250 6.640 2.480 ;
        RECT  2.305 2.780 2.800 3.080 ;
        RECT  2.570 1.915 2.800 3.395 ;
        RECT  2.570 3.165 6.270 3.395 ;
        RECT  5.930 2.250 6.270 3.550 ;
        RECT  7.430 2.075 8.680 2.415 ;
        RECT  7.430 1.240 7.770 3.550 ;
        RECT  0.170 3.380 1.50 3.610 ;
        RECT  2.570 3.165 5.70 3.395 ;
    END
END DLLSQX4

MACRO DLLSQX2
    CLASS CORE ;
    FOREIGN DLLSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 2.640 8.070 3.480 ;
        RECT  7.840 1.240 8.070 3.480 ;
        RECT  7.680 1.240 8.070 1.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.795 2.130 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 1.640 1.135 2.465 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.080 1.585 5.645 2.020 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.920 -0.400 8.580 0.720 ;
        RECT  4.940 -0.400 5.280 1.320 ;
        RECT  3.445 -0.400 3.785 0.955 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.120 4.170 8.580 5.280 ;
        RECT  5.025 3.700 5.365 5.280 ;
        RECT  3.850 3.875 4.190 5.280 ;
        RECT  1.440 4.170 1.780 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.950 ;
        RECT  0.180 0.630 0.410 2.925 ;
        RECT  1.365 1.890 1.650 2.925 ;
        RECT  0.180 2.695 1.650 2.925 ;
        RECT  0.740 2.695 1.080 3.150 ;
        RECT  1.880 1.270 2.585 1.610 ;
        RECT  0.170 3.155 0.510 3.610 ;
        RECT  0.170 3.380 2.110 3.610 ;
        RECT  1.880 1.270 2.110 3.935 ;
        RECT  1.880 3.705 2.960 3.935 ;
        RECT  2.620 3.705 2.960 4.240 ;
        RECT  1.965 0.680 3.045 1.020 ;
        RECT  4.025 0.980 4.560 1.320 ;
        RECT  2.815 0.680 3.045 3.010 ;
        RECT  4.025 0.980 4.255 3.010 ;
        RECT  2.815 2.670 4.255 3.010 ;
        RECT  2.815 2.710 4.605 3.010 ;
        RECT  5.660 0.980 6.125 1.320 ;
        RECT  4.505 2.080 4.845 2.480 ;
        RECT  4.505 2.250 6.125 2.480 ;
        RECT  2.340 2.090 2.585 3.470 ;
        RECT  5.785 2.250 6.125 3.470 ;
        RECT  5.890 0.980 6.125 3.470 ;
        RECT  2.340 3.240 6.125 3.470 ;
        RECT  6.360 1.880 7.610 2.220 ;
        RECT  6.360 1.170 6.700 3.540 ;
        RECT  2.340 3.240 5.70 3.470 ;
    END
END DLLSQX2

MACRO DLLSQX1
    CLASS CORE ;
    FOREIGN DLLSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 3.270 8.695 4.180 ;
        RECT  8.465 0.820 8.695 4.180 ;
        RECT  8.300 0.820 8.695 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.510 4.350 2.220 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.860 1.975 3.270 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.020 6.030 2.360 ;
        RECT  5.165 2.020 5.585 2.630 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.060 ;
        RECT  5.330 -0.400 5.670 1.040 ;
        RECT  3.870 -0.400 4.210 1.280 ;
        RECT  1.210 -0.400 1.550 0.715 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 3.330 7.920 5.280 ;
        RECT  5.400 3.525 5.740 5.280 ;
        RECT  4.290 3.825 4.630 5.280 ;
        RECT  1.655 3.840 1.975 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.120 1.035 0.520 1.465 ;
        RECT  0.120 1.235 1.970 1.465 ;
        RECT  1.630 1.235 1.970 2.170 ;
        RECT  0.120 1.035 0.350 3.250 ;
        RECT  0.120 3.020 1.120 3.250 ;
        RECT  0.890 3.020 1.120 4.175 ;
        RECT  0.890 3.835 1.280 4.175 ;
        RECT  2.205 1.250 2.810 1.590 ;
        RECT  0.580 2.290 0.865 2.630 ;
        RECT  0.580 2.400 2.435 2.630 ;
        RECT  2.205 1.250 2.435 4.115 ;
        RECT  2.205 3.775 3.230 4.115 ;
        RECT  2.190 0.630 3.530 0.970 ;
        RECT  4.580 0.770 4.950 1.120 ;
        RECT  3.300 0.630 3.530 2.835 ;
        RECT  3.300 2.470 3.640 2.835 ;
        RECT  4.580 0.770 4.810 2.835 ;
        RECT  3.300 2.550 4.925 2.835 ;
        RECT  6.045 0.860 6.390 1.790 ;
        RECT  5.055 1.460 6.500 1.790 ;
        RECT  2.665 2.950 2.950 3.295 ;
        RECT  6.150 2.595 6.500 3.295 ;
        RECT  2.665 3.065 6.500 3.295 ;
        RECT  6.260 1.460 6.500 3.350 ;
        RECT  6.160 2.550 6.500 3.350 ;
        RECT  6.780 0.940 7.155 4.180 ;
        RECT  6.780 2.160 8.160 2.500 ;
        RECT  6.780 2.160 7.160 4.180 ;
        RECT  2.665 3.065 5.30 3.295 ;
    END
END DLLSQX1

MACRO DLLSQX0
    CLASS CORE ;
    FOREIGN DLLSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.555 2.995 8.075 3.335 ;
        RECT  7.845 1.260 8.075 3.335 ;
        RECT  7.665 1.260 8.075 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.460 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.760 1.765 3.350 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.930 2.230 5.270 2.755 ;
        RECT  4.535 2.230 5.270 2.630 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.595 -0.400 7.940 0.900 ;
        RECT  5.450 -0.400 6.365 1.145 ;
        RECT  3.950 -0.400 4.290 1.540 ;
        RECT  1.320 -0.400 1.660 1.460 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.055 3.840 7.840 5.280 ;
        RECT  4.450 3.965 5.630 5.280 ;
        RECT  1.755 3.580 2.095 5.280 ;
        RECT  0.180 3.930 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.970 ;
        RECT  0.115 1.740 1.765 1.970 ;
        RECT  1.425 1.740 1.765 2.070 ;
        RECT  0.115 1.740 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  1.995 1.230 2.890 1.540 ;
        RECT  0.575 2.300 2.225 2.530 ;
        RECT  0.575 2.300 0.915 2.955 ;
        RECT  1.995 1.230 2.225 3.240 ;
        RECT  1.995 3.010 3.210 3.240 ;
        RECT  2.980 3.010 3.210 4.250 ;
        RECT  2.980 3.930 3.320 4.250 ;
        RECT  4.560 0.780 4.990 1.120 ;
        RECT  4.650 0.780 4.990 2.000 ;
        RECT  4.650 1.770 5.905 2.000 ;
        RECT  5.600 1.770 5.905 2.365 ;
        RECT  5.600 1.770 5.830 3.275 ;
        RECT  4.690 2.985 5.830 3.275 ;
        RECT  2.455 1.770 2.740 2.580 ;
        RECT  2.455 2.350 3.840 2.580 ;
        RECT  3.445 2.350 3.840 2.635 ;
        RECT  3.445 2.350 3.800 2.655 ;
        RECT  3.445 2.350 3.675 3.735 ;
        RECT  6.080 3.095 6.365 3.735 ;
        RECT  6.135 1.505 6.365 3.735 ;
        RECT  3.445 3.505 6.365 3.735 ;
        RECT  6.595 0.655 7.200 0.995 ;
        RECT  6.595 2.275 7.615 2.615 ;
        RECT  6.595 0.655 6.825 4.250 ;
        RECT  6.180 3.965 6.825 4.250 ;
        RECT  3.445 3.505 5.20 3.735 ;
    END
END DLLSQX0

MACRO DLLRX4
    CLASS CORE ;
    FOREIGN DLLRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 1.240 13.105 4.100 ;
        RECT  11.550 2.250 13.105 2.480 ;
        RECT  11.390 2.640 11.780 3.770 ;
        RECT  11.550 0.790 11.780 3.770 ;
        RECT  11.390 0.790 11.780 1.700 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.900 3.025 6.280 3.385 ;
        RECT  5.780 2.855 6.240 3.260 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.550 1.135 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.070 1.240 10.410 3.450 ;
        RECT  8.750 2.250 10.410 2.630 ;
        RECT  8.750 1.240 9.090 3.450 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  12.150 -0.400 12.490 0.720 ;
        RECT  6.870 -0.400 10.970 0.720 ;
        RECT  5.450 -0.400 5.790 1.205 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  7.990 4.140 12.290 5.280 ;
        RECT  6.670 2.925 7.010 5.280 ;
        RECT  4.545 4.150 4.885 5.280 ;
        RECT  2.205 3.900 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  1.350 2.105 1.670 2.480 ;
        RECT  1.360 2.080 1.670 2.480 ;
        RECT  0.180 2.250 1.670 2.480 ;
        RECT  3.875 2.455 4.215 2.795 ;
        RECT  0.180 2.250 0.520 3.460 ;
        RECT  3.875 2.455 4.105 3.460 ;
        RECT  0.180 3.230 4.105 3.460 ;
        RECT  1.700 0.980 2.130 1.320 ;
        RECT  3.940 1.785 4.225 2.125 ;
        RECT  3.315 1.895 4.225 2.125 ;
        RECT  1.740 2.700 2.130 3.000 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.710 2.130 3.000 ;
        RECT  3.155 2.700 3.545 3.000 ;
        RECT  3.315 1.895 3.545 3.000 ;
        RECT  1.700 2.770 3.545 3.000 ;
        RECT  2.460 0.630 5.145 0.955 ;
        RECT  4.915 0.630 5.145 1.665 ;
        RECT  6.170 0.950 6.510 1.665 ;
        RECT  4.915 1.435 6.510 1.665 ;
        RECT  3.660 1.215 4.000 1.555 ;
        RECT  3.660 1.325 4.685 1.555 ;
        RECT  4.455 1.895 7.200 2.125 ;
        RECT  6.860 1.895 7.200 2.235 ;
        RECT  4.455 1.325 4.685 3.920 ;
        RECT  4.455 3.580 5.685 3.920 ;
        RECT  3.435 3.690 5.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  10.785 2.075 11.320 2.415 ;
        RECT  4.915 2.355 6.630 2.585 ;
        RECT  4.915 2.355 5.200 2.695 ;
        RECT  6.410 2.465 7.770 2.695 ;
        RECT  7.430 1.240 7.770 3.910 ;
        RECT  10.785 2.075 11.015 3.910 ;
        RECT  7.430 3.680 11.015 3.910 ;
        RECT  0.180 3.230 3.60 3.460 ;
        RECT  2.460 0.630 4.80 0.955 ;
        RECT  4.455 1.895 6.90 2.125 ;
        RECT  3.435 3.690 4.50 3.920 ;
        RECT  7.430 3.680 10.60 3.910 ;
    END
END DLLRX4

MACRO DLLRX2
    CLASS CORE ;
    FOREIGN DLLRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.240 1.135 3.480 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.400 2.595 4.915 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.015 1.640 7.575 2.085 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 1.550 9.435 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.240 2.400 3.480 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.800 -0.400 9.140 1.320 ;
        RECT  0.180 -0.400 4.220 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.800 3.685 9.140 5.280 ;
        RECT  7.485 3.685 7.825 5.280 ;
        RECT  5.195 3.930 5.535 5.280 ;
        RECT  1.500 4.170 2.960 5.280 ;
        RECT  0.180 4.010 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.270 1.240 3.720 1.795 ;
        RECT  3.270 1.565 5.115 1.795 ;
        RECT  4.830 1.565 5.115 1.905 ;
        RECT  3.270 2.640 3.720 3.550 ;
        RECT  3.270 1.240 3.500 3.940 ;
        RECT  0.930 3.710 3.500 3.940 ;
        RECT  0.930 3.710 1.270 4.070 ;
        RECT  5.345 1.090 6.210 1.335 ;
        RECT  3.730 2.025 4.070 2.365 ;
        RECT  3.730 2.135 5.575 2.365 ;
        RECT  5.345 1.090 5.575 3.700 ;
        RECT  4.395 3.470 6.595 3.700 ;
        RECT  4.395 3.470 4.735 3.810 ;
        RECT  6.255 3.470 6.595 3.810 ;
        RECT  4.640 0.630 7.640 0.860 ;
        RECT  4.640 0.630 4.980 1.215 ;
        RECT  7.300 0.630 7.640 1.310 ;
        RECT  7.950 0.980 8.380 1.320 ;
        RECT  5.805 1.565 6.090 1.905 ;
        RECT  5.805 1.675 6.765 1.905 ;
        RECT  6.535 1.675 6.765 2.780 ;
        RECT  6.535 2.480 6.875 2.780 ;
        RECT  7.950 0.980 8.180 2.995 ;
        RECT  6.535 2.700 8.340 2.780 ;
        RECT  6.535 2.550 8.180 2.780 ;
        RECT  7.950 2.710 8.380 2.995 ;
        RECT  9.560 0.980 9.900 1.320 ;
        RECT  8.410 2.080 8.720 2.480 ;
        RECT  8.410 2.105 8.730 2.480 ;
        RECT  8.410 2.250 9.900 2.480 ;
        RECT  5.865 2.235 6.205 2.575 ;
        RECT  5.975 2.235 6.205 3.240 ;
        RECT  9.560 2.250 9.900 3.455 ;
        RECT  5.975 3.010 7.405 3.240 ;
        RECT  9.665 0.980 9.900 3.455 ;
        RECT  7.175 3.225 9.900 3.455 ;
        RECT  0.930 3.710 2.70 3.940 ;
        RECT  4.395 3.470 5.60 3.700 ;
        RECT  4.640 0.630 6.90 0.860 ;
        RECT  7.175 3.225 8.70 3.455 ;
    END
END DLLRX2

MACRO DLLRX1
    CLASS CORE ;
    FOREIGN DLLRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.820 0.520 3.880 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.110 1.615 3.665 2.060 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 2.970 1.960 3.780 ;
        RECT  1.620 0.700 1.960 1.040 ;
        RECT  1.620 0.700 1.850 1.495 ;
        RECT  1.385 2.250 1.765 2.630 ;
        RECT  1.470 1.265 1.700 3.215 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.470 2.095 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.975 8.160 2.315 ;
        RECT  7.685 1.975 8.145 2.635 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.575 -0.400 7.915 1.270 ;
        RECT  2.765 -0.400 3.105 0.710 ;
        RECT  0.900 -0.400 1.240 1.060 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.540 3.525 7.880 5.280 ;
        RECT  6.440 3.800 6.780 5.280 ;
        RECT  3.095 3.530 4.130 5.280 ;
        RECT  0.900 3.030 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.160 1.360 2.500 1.700 ;
        RECT  2.160 1.360 2.425 2.350 ;
        RECT  1.995 2.010 2.425 2.350 ;
        RECT  2.195 1.360 2.425 3.850 ;
        RECT  2.195 3.510 2.715 3.850 ;
        RECT  4.755 1.090 5.095 1.375 ;
        RECT  4.070 1.145 5.095 1.375 ;
        RECT  2.655 2.440 2.955 3.050 ;
        RECT  4.070 1.145 4.300 3.050 ;
        RECT  2.655 2.710 4.300 3.050 ;
        RECT  2.655 2.750 4.590 3.050 ;
        RECT  4.360 2.750 4.590 3.940 ;
        RECT  4.360 3.600 5.420 3.940 ;
        RECT  3.525 0.630 6.495 0.860 ;
        RECT  3.525 0.630 3.865 1.040 ;
        RECT  6.155 0.630 6.495 1.375 ;
        RECT  6.855 0.810 7.195 1.730 ;
        RECT  4.530 1.605 5.545 1.945 ;
        RECT  5.315 1.605 5.545 2.835 ;
        RECT  5.315 2.415 5.830 2.835 ;
        RECT  6.740 1.495 6.970 2.835 ;
        RECT  5.315 2.550 6.970 2.835 ;
        RECT  8.295 0.865 8.640 1.205 ;
        RECT  7.200 1.980 7.455 3.295 ;
        RECT  8.290 2.820 8.640 3.295 ;
        RECT  8.405 0.865 8.640 3.295 ;
        RECT  4.820 3.065 8.640 3.295 ;
        RECT  4.820 3.010 5.160 3.350 ;
        RECT  3.525 0.630 5.60 0.860 ;
        RECT  4.820 3.065 7.70 3.295 ;
    END
END DLLRX1

MACRO DLLRX0
    CLASS CORE ;
    FOREIGN DLLRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.910 2.250 5.545 2.630 ;
        RECT  4.910 1.890 5.250 2.630 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.469  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.925 3.130 7.445 3.470 ;
        RECT  7.215 0.630 7.445 3.470 ;
        RECT  7.055 2.250 7.445 2.630 ;
        RECT  6.690 0.630 7.445 0.960 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.443  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.880 6.175 3.170 ;
        RECT  5.775 1.030 6.175 1.410 ;
        RECT  5.775 1.030 6.005 3.170 ;
        RECT  5.260 1.250 6.005 1.605 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.180 2.595 2.630 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 2.190 1.765 2.630 ;
        END
    END GN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.925 3.930 7.265 5.280 ;
        RECT  4.110 3.860 5.330 5.280 ;
        RECT  0.880 3.895 1.820 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.210 -0.400 6.205 0.800 ;
        RECT  0.880 -0.400 1.220 1.060 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.480 0.630 1.820 1.700 ;
        RECT  0.750 1.470 1.820 1.700 ;
        RECT  0.575 1.935 0.980 2.275 ;
        RECT  0.750 1.470 0.980 3.090 ;
        RECT  0.750 2.860 1.820 3.090 ;
        RECT  1.480 2.860 1.820 3.205 ;
        RECT  0.115 0.720 0.520 1.060 ;
        RECT  3.625 1.915 3.965 2.255 ;
        RECT  3.625 1.915 3.855 3.090 ;
        RECT  2.420 2.860 3.855 3.090 ;
        RECT  2.420 2.860 2.770 3.190 ;
        RECT  0.115 0.720 0.345 3.995 ;
        RECT  2.420 2.860 2.650 3.665 ;
        RECT  0.115 3.435 2.650 3.665 ;
        RECT  0.115 3.435 0.520 3.995 ;
        RECT  2.180 0.680 4.750 0.910 ;
        RECT  2.180 0.680 2.520 1.020 ;
        RECT  4.410 0.680 4.750 1.035 ;
        RECT  3.380 1.195 3.720 1.535 ;
        RECT  3.380 1.305 4.540 1.535 ;
        RECT  4.310 1.305 4.540 3.630 ;
        RECT  4.310 2.985 4.730 3.630 ;
        RECT  2.880 3.400 6.235 3.630 ;
        RECT  5.910 3.400 6.235 3.750 ;
        RECT  2.880 3.400 3.220 3.885 ;
        RECT  6.465 1.320 6.985 1.660 ;
        RECT  6.235 2.305 6.695 2.645 ;
        RECT  6.465 1.320 6.695 4.250 ;
        RECT  6.035 3.980 6.695 4.250 ;
        RECT  0.115 3.435 1.60 3.665 ;
        RECT  2.180 0.680 3.80 0.910 ;
        RECT  2.880 3.400 5.30 3.630 ;
    END
END DLLRX0

MACRO DLLRSX4
    CLASS CORE ;
    FOREIGN DLLRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.875 1.550 7.435 2.020 ;
        END
    END GN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.330 1.240 11.670 3.450 ;
        RECT  10.010 2.250 11.670 2.630 ;
        RECT  10.010 1.240 10.350 3.450 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.140 2.030 2.480 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.140 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.065 1.640 5.545 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 1.240 14.365 4.100 ;
        RECT  12.810 2.250 14.365 2.480 ;
        RECT  12.650 2.640 13.040 3.770 ;
        RECT  12.810 0.790 13.040 3.770 ;
        RECT  12.650 0.790 13.040 1.700 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.410 -0.400 13.750 0.720 ;
        RECT  8.130 -0.400 12.230 0.720 ;
        RECT  6.710 -0.400 7.050 1.320 ;
        RECT  2.330 -0.400 2.670 0.655 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  9.250 4.140 13.550 5.280 ;
        RECT  7.970 2.710 8.310 5.280 ;
        RECT  6.430 3.625 6.770 5.280 ;
        RECT  5.185 3.900 5.525 5.280 ;
        RECT  1.540 3.930 2.920 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.910 ;
        RECT  1.365 1.680 2.730 1.910 ;
        RECT  2.500 1.680 2.730 2.610 ;
        RECT  2.510 2.290 2.840 2.625 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  4.060 1.235 4.400 1.575 ;
        RECT  3.070 1.345 4.400 1.575 ;
        RECT  1.995 2.740 2.310 3.700 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.995 2.775 2.335 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 3.525 3.700 ;
        RECT  3.070 1.345 3.300 3.700 ;
        RECT  3.300 3.625 4.225 3.855 ;
        RECT  3.885 3.625 4.225 3.965 ;
        RECT  3.030 0.670 5.630 0.970 ;
        RECT  5.290 0.630 5.630 0.970 ;
        RECT  1.825 0.885 3.370 1.115 ;
        RECT  1.825 0.885 2.110 1.450 ;
        RECT  5.990 0.980 6.330 1.385 ;
        RECT  5.780 1.155 6.010 2.935 ;
        RECT  4.235 2.595 6.010 2.935 ;
        RECT  7.430 0.980 7.900 1.320 ;
        RECT  3.775 1.805 4.835 2.145 ;
        RECT  6.240 2.120 6.570 2.480 ;
        RECT  7.665 0.980 7.900 2.480 ;
        RECT  6.240 2.250 7.900 2.480 ;
        RECT  3.530 2.740 4.005 3.080 ;
        RECT  3.775 1.805 4.005 3.395 ;
        RECT  3.775 3.165 7.530 3.395 ;
        RECT  7.190 2.250 7.530 3.550 ;
        RECT  12.190 2.075 12.580 2.415 ;
        RECT  8.690 1.240 9.030 3.910 ;
        RECT  12.190 2.075 12.420 3.910 ;
        RECT  8.690 3.680 12.420 3.910 ;
        RECT  0.965 3.470 2.40 3.700 ;
        RECT  3.030 0.670 4.60 0.970 ;
        RECT  3.775 3.165 6.70 3.395 ;
        RECT  8.690 3.680 11.60 3.910 ;
    END
END DLLRSX4

MACRO DLLRSX2
    CLASS CORE ;
    FOREIGN DLLRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.940 1.240 9.325 3.480 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.280 2.030 2.620 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.280 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.500 1.640 5.055 2.080 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.075 1.200 2.410 ;
        RECT  0.755 1.640 1.135 2.410 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 1.240 10.600 3.480 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.345 1.560 6.905 2.020 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  8.180 -0.400 11.160 0.720 ;
        RECT  6.045 -0.400 6.385 1.320 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 4.010 11.160 5.280 ;
        RECT  8.380 4.170 9.840 5.280 ;
        RECT  6.285 3.630 6.625 5.280 ;
        RECT  4.970 3.630 5.310 5.280 ;
        RECT  1.540 3.930 2.900 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.795 ;
        RECT  1.365 1.565 2.245 1.795 ;
        RECT  1.960 1.565 2.245 1.905 ;
        RECT  0.180 0.630 0.410 2.870 ;
        RECT  0.180 2.640 1.080 2.870 ;
        RECT  0.740 2.640 1.080 3.150 ;
        RECT  2.475 1.090 3.340 1.335 ;
        RECT  0.170 3.100 0.510 3.610 ;
        RECT  2.475 1.090 2.705 3.700 ;
        RECT  1.995 2.850 2.705 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 4.080 3.700 ;
        RECT  3.740 3.470 4.080 4.010 ;
        RECT  1.775 0.630 4.770 0.860 ;
        RECT  1.775 0.630 2.110 1.035 ;
        RECT  1.785 0.630 2.110 1.045 ;
        RECT  4.430 0.630 4.770 1.310 ;
        RECT  5.285 0.980 5.625 1.320 ;
        RECT  2.935 1.565 3.220 1.905 ;
        RECT  2.935 1.675 4.250 1.905 ;
        RECT  4.020 1.675 4.250 2.630 ;
        RECT  4.020 2.290 4.360 2.630 ;
        RECT  4.020 2.400 5.515 2.630 ;
        RECT  5.285 0.980 5.515 2.940 ;
        RECT  5.285 2.710 5.865 2.940 ;
        RECT  6.805 0.980 7.385 1.320 ;
        RECT  5.765 2.080 6.105 2.480 ;
        RECT  5.765 2.250 7.385 2.480 ;
        RECT  3.350 2.180 3.690 2.520 ;
        RECT  3.460 2.180 3.690 3.240 ;
        RECT  7.045 2.250 7.385 3.400 ;
        RECT  3.460 3.010 4.890 3.240 ;
        RECT  7.150 0.980 7.385 3.400 ;
        RECT  4.660 3.170 7.385 3.400 ;
        RECT  7.620 1.170 7.960 3.940 ;
        RECT  7.620 3.710 10.410 3.940 ;
        RECT  10.070 3.710 10.410 4.070 ;
        RECT  0.965 3.470 3.60 3.700 ;
        RECT  1.775 0.630 3.90 0.860 ;
        RECT  4.660 3.170 6.70 3.400 ;
        RECT  7.620 3.710 9.00 3.940 ;
    END
END DLLRSX2

MACRO DLLRSX1
    CLASS CORE ;
    FOREIGN DLLRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.860 2.250 9.325 2.630 ;
        RECT  8.750 3.270 9.090 4.080 ;
        RECT  8.860 0.700 9.090 4.080 ;
        RECT  8.750 0.700 9.090 1.040 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.810 2.230 2.400 2.665 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 0.820 10.585 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.285 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.400 2.070 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.665 1.500 7.005 1.840 ;
        RECT  6.665 1.030 6.955 1.840 ;
        RECT  6.425 1.030 6.955 1.415 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.060 ;
        RECT  7.950 -0.400 8.290 0.710 ;
        RECT  6.295 -0.400 6.635 0.710 ;
        RECT  1.210 -0.400 1.550 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 3.330 9.810 5.280 ;
        RECT  7.815 4.170 8.155 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.630 0.520 1.410 ;
        RECT  0.170 1.210 1.860 1.410 ;
        RECT  0.170 1.180 1.835 1.410 ;
        RECT  1.630 1.335 2.445 1.680 ;
        RECT  0.170 0.630 0.400 3.250 ;
        RECT  0.170 3.020 1.120 3.250 ;
        RECT  0.780 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 1.580 2.785 ;
        RECT  1.350 2.445 1.580 3.340 ;
        RECT  1.350 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  2.000 0.630 5.135 0.860 ;
        RECT  2.000 0.630 2.310 1.015 ;
        RECT  2.025 0.630 2.310 1.040 ;
        RECT  4.795 0.630 5.135 1.280 ;
        RECT  5.515 0.810 5.875 1.150 ;
        RECT  3.135 1.555 4.305 1.785 ;
        RECT  3.135 1.555 3.420 1.895 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 5.745 2.655 ;
        RECT  5.515 0.810 5.745 2.655 ;
        RECT  5.535 2.550 6.040 2.835 ;
        RECT  7.230 0.980 7.615 1.320 ;
        RECT  5.975 1.760 6.260 2.320 ;
        RECT  5.975 2.075 7.615 2.320 ;
        RECT  3.520 2.500 3.845 3.115 ;
        RECT  7.265 2.720 7.615 3.295 ;
        RECT  3.520 2.885 5.120 3.115 ;
        RECT  7.380 0.980 7.615 3.295 ;
        RECT  4.890 3.065 7.615 3.295 ;
        RECT  7.930 1.170 8.380 1.510 ;
        RECT  7.930 2.130 8.615 2.505 ;
        RECT  7.930 1.170 8.160 3.820 ;
        RECT  7.815 3.445 8.160 3.820 ;
        RECT  2.000 0.630 4.30 0.860 ;
        RECT  4.890 3.065 6.20 3.295 ;
    END
END DLLRSX1

MACRO DLLRSX0
    CLASS CORE ;
    FOREIGN DLLRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.225 2.250 8.065 2.630 ;
        RECT  7.225 0.675 7.870 1.015 ;
        RECT  6.810 3.965 7.455 4.250 ;
        RECT  7.225 0.675 7.455 4.250 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.395 2.630 ;
        RECT  1.790 2.120 2.395 2.460 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.578  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 0.630 9.335 4.135 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.090 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.270 2.280 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.560 2.230 5.900 2.755 ;
        RECT  5.165 2.230 5.900 2.630 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.225 -0.400 8.570 0.970 ;
        RECT  6.080 -0.400 6.995 1.145 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.685 3.885 8.495 5.280 ;
        RECT  5.190 3.965 6.260 5.280 ;
        RECT  1.645 3.660 2.790 5.280 ;
        RECT  0.180 3.700 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 2.395 1.410 ;
        RECT  2.055 1.180 2.395 1.790 ;
        RECT  0.115 1.200 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  0.900 3.185 1.155 4.000 ;
        RECT  0.900 3.660 1.240 4.000 ;
        RECT  2.625 1.230 3.520 1.540 ;
        RECT  0.575 2.610 0.915 2.955 ;
        RECT  0.575 2.695 1.615 2.955 ;
        RECT  2.625 1.230 2.855 3.200 ;
        RECT  1.385 2.860 2.855 3.200 ;
        RECT  1.385 2.970 3.440 3.200 ;
        RECT  3.210 2.970 3.440 4.250 ;
        RECT  3.210 3.965 4.185 4.250 ;
        RECT  1.950 0.630 2.290 0.950 ;
        RECT  1.950 0.720 4.920 0.950 ;
        RECT  4.580 0.720 4.920 1.540 ;
        RECT  5.180 0.780 5.620 1.120 ;
        RECT  5.280 0.780 5.620 2.000 ;
        RECT  5.280 1.770 6.535 2.000 ;
        RECT  6.230 1.770 6.535 2.365 ;
        RECT  6.230 1.770 6.460 3.275 ;
        RECT  5.320 2.985 6.460 3.275 ;
        RECT  3.085 1.770 3.370 2.580 ;
        RECT  3.085 2.350 4.470 2.580 ;
        RECT  4.075 2.350 4.470 2.635 ;
        RECT  4.075 2.350 4.430 2.655 ;
        RECT  4.075 2.350 4.305 3.735 ;
        RECT  6.710 3.095 6.995 3.735 ;
        RECT  6.765 1.505 6.995 3.735 ;
        RECT  4.075 3.505 6.995 3.735 ;
        RECT  7.685 1.375 8.525 1.715 ;
        RECT  8.295 2.395 8.700 2.735 ;
        RECT  8.295 1.375 8.525 3.420 ;
        RECT  7.745 3.080 8.525 3.420 ;
        RECT  0.180 1.180 1.70 1.410 ;
        RECT  1.385 2.970 2.70 3.200 ;
        RECT  1.950 0.720 3.60 0.950 ;
        RECT  4.075 3.505 5.50 3.735 ;
    END
END DLLRSX0

MACRO DLLRSQX4
    CLASS CORE ;
    FOREIGN DLLRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.840 1.610 7.435 2.020 ;
        END
    END GN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.140 2.030 2.480 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.140 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.065 1.640 5.545 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.450 1.130 11.845 3.880 ;
        RECT  10.170 2.130 11.845 2.360 ;
        RECT  10.010 2.640 10.400 3.880 ;
        RECT  10.170 1.130 10.400 3.880 ;
        RECT  10.010 1.130 10.400 1.470 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.730 -0.400 11.070 1.470 ;
        RECT  8.130 -0.400 9.590 0.720 ;
        RECT  6.710 -0.400 7.050 1.380 ;
        RECT  2.330 -0.400 2.670 0.655 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.730 2.640 11.070 5.280 ;
        RECT  9.250 3.950 9.590 5.280 ;
        RECT  7.970 2.700 8.310 5.280 ;
        RECT  6.430 3.625 6.770 5.280 ;
        RECT  5.185 3.900 5.525 5.280 ;
        RECT  1.540 3.930 2.920 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.910 ;
        RECT  1.365 1.680 2.840 1.910 ;
        RECT  2.500 1.680 2.840 2.610 ;
        RECT  2.510 1.680 2.840 2.625 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  4.060 1.235 4.400 1.575 ;
        RECT  3.070 1.345 4.400 1.575 ;
        RECT  1.995 2.740 2.310 3.700 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.995 2.775 2.335 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 3.525 3.700 ;
        RECT  3.070 1.345 3.300 3.700 ;
        RECT  3.300 3.625 4.225 3.855 ;
        RECT  3.885 3.625 4.225 3.965 ;
        RECT  3.030 0.670 5.630 0.970 ;
        RECT  5.290 0.630 5.630 0.970 ;
        RECT  1.825 0.885 3.370 1.115 ;
        RECT  1.825 0.885 2.110 1.450 ;
        RECT  5.990 1.040 6.330 1.380 ;
        RECT  5.780 1.150 6.010 2.935 ;
        RECT  4.235 2.595 6.010 2.935 ;
        RECT  7.430 1.040 7.900 1.380 ;
        RECT  4.495 1.805 4.835 2.145 ;
        RECT  3.775 1.915 4.835 2.145 ;
        RECT  6.240 2.120 6.570 2.480 ;
        RECT  7.665 1.040 7.900 2.480 ;
        RECT  6.240 2.250 7.900 2.480 ;
        RECT  3.530 2.740 4.005 3.080 ;
        RECT  3.775 1.915 4.005 3.395 ;
        RECT  3.775 3.165 7.530 3.395 ;
        RECT  7.190 2.250 7.530 3.550 ;
        RECT  8.690 2.075 9.940 2.415 ;
        RECT  8.690 1.240 9.030 3.550 ;
        RECT  0.965 3.470 2.80 3.700 ;
        RECT  3.030 0.670 4.20 0.970 ;
        RECT  3.775 3.165 6.30 3.395 ;
    END
END DLLRSQX4

MACRO DLLRSQX2
    CLASS CORE ;
    FOREIGN DLLRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.280 2.030 2.620 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.280 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.500 1.640 5.055 2.080 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.075 1.200 2.410 ;
        RECT  0.755 1.640 1.135 2.410 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.375 1.570 6.920 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.640 9.390 3.550 ;
        RECT  9.160 1.240 9.390 3.550 ;
        RECT  9.000 1.240 9.390 1.580 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.240 -0.400 9.900 0.720 ;
        RECT  6.045 -0.400 6.385 1.320 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.440 3.950 9.900 5.280 ;
        RECT  6.285 3.630 6.625 5.280 ;
        RECT  4.970 3.630 5.310 5.280 ;
        RECT  1.540 3.930 2.900 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.795 ;
        RECT  1.365 1.565 2.245 1.795 ;
        RECT  1.960 1.565 2.245 1.905 ;
        RECT  0.180 0.630 0.410 2.870 ;
        RECT  0.180 2.640 1.080 2.870 ;
        RECT  0.740 2.640 1.080 3.150 ;
        RECT  2.475 1.090 3.340 1.335 ;
        RECT  0.170 3.100 0.510 3.610 ;
        RECT  2.475 1.090 2.705 3.700 ;
        RECT  1.995 2.850 2.705 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 4.080 3.700 ;
        RECT  3.740 3.470 4.080 4.010 ;
        RECT  1.775 0.630 4.770 0.860 ;
        RECT  1.775 0.630 2.110 1.035 ;
        RECT  1.785 0.630 2.110 1.045 ;
        RECT  4.430 0.630 4.770 1.310 ;
        RECT  5.285 0.980 5.625 1.320 ;
        RECT  2.935 1.565 3.220 1.905 ;
        RECT  2.935 1.675 4.250 1.905 ;
        RECT  4.020 1.675 4.250 2.630 ;
        RECT  4.020 2.290 4.360 2.630 ;
        RECT  4.020 2.400 5.515 2.630 ;
        RECT  5.285 0.980 5.515 2.940 ;
        RECT  5.285 2.710 5.865 2.940 ;
        RECT  6.805 0.980 7.385 1.320 ;
        RECT  5.765 2.080 6.105 2.480 ;
        RECT  5.765 2.250 7.385 2.480 ;
        RECT  3.350 2.180 3.690 2.520 ;
        RECT  3.460 2.180 3.690 3.240 ;
        RECT  7.045 2.250 7.385 3.400 ;
        RECT  3.460 3.010 4.890 3.240 ;
        RECT  7.150 0.980 7.385 3.400 ;
        RECT  4.660 3.170 7.385 3.400 ;
        RECT  7.680 2.040 8.930 2.270 ;
        RECT  8.590 2.040 8.930 2.380 ;
        RECT  7.680 1.240 8.020 3.550 ;
        RECT  0.965 3.470 3.20 3.700 ;
        RECT  1.775 0.630 3.50 0.860 ;
        RECT  4.660 3.170 6.10 3.400 ;
    END
END DLLRSQX2

MACRO DLLRSQX1
    CLASS CORE ;
    FOREIGN DLLRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.810 2.230 2.400 2.665 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.560 0.820 9.955 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.285 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.400 2.070 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.665 1.030 7.005 1.840 ;
        RECT  6.425 1.030 7.005 1.415 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.840 -0.400 9.180 1.140 ;
        RECT  6.295 -0.400 6.635 0.710 ;
        RECT  1.210 -0.400 1.550 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.840 3.330 9.180 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.630 0.520 1.410 ;
        RECT  0.170 1.210 1.860 1.410 ;
        RECT  0.170 1.180 1.835 1.410 ;
        RECT  1.630 1.335 2.445 1.680 ;
        RECT  0.170 0.630 0.400 3.360 ;
        RECT  0.170 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 1.580 2.785 ;
        RECT  1.350 2.445 1.580 3.340 ;
        RECT  1.350 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  1.995 0.630 5.025 0.860 ;
        RECT  4.795 0.630 5.025 1.280 ;
        RECT  1.995 0.630 2.310 1.010 ;
        RECT  2.025 0.630 2.310 1.040 ;
        RECT  4.795 0.940 5.135 1.280 ;
        RECT  5.515 0.810 5.875 1.150 ;
        RECT  3.135 1.555 4.305 1.895 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 5.745 2.655 ;
        RECT  5.515 0.810 5.745 2.655 ;
        RECT  5.535 2.550 6.040 2.835 ;
        RECT  5.995 1.980 6.335 2.320 ;
        RECT  5.995 2.075 7.615 2.320 ;
        RECT  3.520 2.500 3.845 3.115 ;
        RECT  3.520 2.885 5.120 3.115 ;
        RECT  7.235 0.835 7.615 3.295 ;
        RECT  4.890 3.065 7.615 3.295 ;
        RECT  8.040 2.160 8.635 2.500 ;
        RECT  8.040 0.700 8.425 3.610 ;
        RECT  1.995 0.630 4.40 0.860 ;
        RECT  4.890 3.065 6.80 3.295 ;
    END
END DLLRSQX1

MACRO DLLRSQX0
    CLASS CORE ;
    FOREIGN DLLRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.395 2.630 ;
        RECT  1.790 2.120 2.395 2.460 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.185 2.995 8.705 3.335 ;
        RECT  8.475 1.260 8.705 3.335 ;
        RECT  8.295 1.260 8.705 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.090 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.270 2.280 ;
        END
    END SN
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.560 2.230 5.900 2.755 ;
        RECT  5.165 2.230 5.900 2.630 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.225 -0.400 8.570 0.900 ;
        RECT  6.080 -0.400 6.995 1.145 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.685 3.795 8.470 5.280 ;
        RECT  5.080 3.965 6.260 5.280 ;
        RECT  1.645 3.660 2.865 5.280 ;
        RECT  0.180 3.700 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.410 ;
        RECT  0.115 1.180 2.395 1.410 ;
        RECT  2.055 1.180 2.395 1.790 ;
        RECT  0.115 0.630 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  0.900 3.185 1.155 4.000 ;
        RECT  0.900 3.660 1.240 4.000 ;
        RECT  2.625 1.230 3.520 1.540 ;
        RECT  0.575 2.610 0.915 2.955 ;
        RECT  0.575 2.695 1.615 2.955 ;
        RECT  2.625 1.230 2.855 3.200 ;
        RECT  1.385 2.860 2.855 3.200 ;
        RECT  1.385 2.970 3.840 3.200 ;
        RECT  3.610 2.970 3.840 4.250 ;
        RECT  3.610 3.965 4.185 4.250 ;
        RECT  1.950 0.630 4.920 0.950 ;
        RECT  4.580 0.630 4.920 1.645 ;
        RECT  5.180 0.780 5.620 1.120 ;
        RECT  5.280 0.780 5.620 2.000 ;
        RECT  5.280 1.770 6.535 2.000 ;
        RECT  6.230 1.770 6.535 2.365 ;
        RECT  6.230 1.770 6.460 3.275 ;
        RECT  5.320 2.985 6.460 3.275 ;
        RECT  3.085 1.770 3.370 2.580 ;
        RECT  3.085 2.350 4.470 2.580 ;
        RECT  4.075 2.350 4.470 2.635 ;
        RECT  4.075 2.350 4.430 2.655 ;
        RECT  4.075 2.350 4.305 3.735 ;
        RECT  6.710 3.095 6.995 3.735 ;
        RECT  6.765 1.505 6.995 3.735 ;
        RECT  4.075 3.505 6.995 3.735 ;
        RECT  7.225 0.655 7.850 0.995 ;
        RECT  7.225 2.275 8.155 2.615 ;
        RECT  7.225 0.655 7.455 4.250 ;
        RECT  6.810 3.965 7.455 4.250 ;
        RECT  0.115 1.180 1.40 1.410 ;
        RECT  1.385 2.970 2.40 3.200 ;
        RECT  1.950 0.630 3.30 0.950 ;
        RECT  4.075 3.505 5.20 3.735 ;
    END
END DLLRSQX0

MACRO DLLRQX4
    CLASS CORE ;
    FOREIGN DLLRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.900 3.025 6.280 3.385 ;
        RECT  5.780 2.855 6.240 3.260 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.550 1.135 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 1.130 10.585 3.880 ;
        RECT  8.750 2.180 10.585 2.410 ;
        RECT  8.750 1.130 9.090 3.880 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.470 ;
        RECT  6.870 -0.400 8.330 0.720 ;
        RECT  5.450 -0.400 5.790 1.205 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 2.640 9.810 5.280 ;
        RECT  7.990 4.140 8.330 5.280 ;
        RECT  6.670 2.925 7.010 5.280 ;
        RECT  4.545 4.150 4.885 5.280 ;
        RECT  2.205 3.900 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  1.350 2.105 1.670 2.480 ;
        RECT  1.360 2.080 1.670 2.480 ;
        RECT  0.180 2.250 1.670 2.480 ;
        RECT  0.180 2.250 0.520 3.460 ;
        RECT  3.875 2.455 4.215 3.460 ;
        RECT  0.180 3.230 4.215 3.460 ;
        RECT  1.700 0.980 2.130 1.320 ;
        RECT  3.315 1.785 4.225 2.125 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.740 2.700 3.545 3.000 ;
        RECT  3.315 1.785 3.545 3.000 ;
        RECT  1.700 2.710 3.545 3.000 ;
        RECT  2.460 0.630 5.145 0.955 ;
        RECT  4.915 0.630 5.145 1.665 ;
        RECT  6.170 0.950 6.510 1.665 ;
        RECT  4.915 1.435 6.510 1.665 ;
        RECT  3.660 1.215 4.685 1.555 ;
        RECT  4.455 1.895 7.200 2.125 ;
        RECT  6.860 1.895 7.200 2.235 ;
        RECT  4.455 1.215 4.685 3.920 ;
        RECT  4.455 3.580 5.685 3.920 ;
        RECT  3.435 3.690 5.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  4.915 2.355 6.630 2.585 ;
        RECT  4.915 2.355 5.200 2.695 ;
        RECT  6.410 2.465 7.770 2.695 ;
        RECT  7.430 1.240 7.770 3.550 ;
        RECT  0.180 3.230 3.50 3.460 ;
        RECT  2.460 0.630 4.00 0.955 ;
        RECT  4.455 1.895 6.40 2.125 ;
        RECT  3.435 3.690 4.80 3.920 ;
    END
END DLLRQX4

MACRO DLLRQX2
    CLASS CORE ;
    FOREIGN DLLRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.550 8.175 2.020 ;
        END
    END GN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.140 2.595 3.655 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.755 1.640 6.315 2.085 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.240 1.140 3.480 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.540 -0.400 7.880 1.320 ;
        RECT  0.240 -0.400 2.960 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.540 3.740 7.880 5.280 ;
        RECT  6.225 3.740 6.565 5.280 ;
        RECT  3.935 3.930 4.275 5.280 ;
        RECT  0.240 4.170 1.700 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.010 1.240 2.460 1.795 ;
        RECT  2.010 1.565 3.855 1.795 ;
        RECT  3.570 1.565 3.855 1.905 ;
        RECT  2.010 1.240 2.240 3.550 ;
        RECT  2.010 2.640 2.460 3.550 ;
        RECT  4.085 1.090 4.950 1.335 ;
        RECT  2.470 2.025 2.810 2.365 ;
        RECT  2.470 2.135 4.315 2.365 ;
        RECT  4.085 1.090 4.315 3.700 ;
        RECT  3.135 3.470 5.335 3.700 ;
        RECT  3.135 3.470 3.475 3.810 ;
        RECT  4.995 3.470 5.335 3.810 ;
        RECT  3.380 0.630 6.270 0.860 ;
        RECT  6.040 0.630 6.270 1.310 ;
        RECT  3.380 0.630 3.720 1.215 ;
        RECT  6.040 0.970 6.380 1.310 ;
        RECT  6.690 0.980 7.120 1.320 ;
        RECT  4.545 1.565 5.505 1.905 ;
        RECT  5.275 1.565 5.505 2.780 ;
        RECT  6.690 0.980 6.920 3.050 ;
        RECT  5.275 2.480 6.920 2.780 ;
        RECT  6.690 2.710 7.120 3.050 ;
        RECT  8.300 0.980 8.640 1.320 ;
        RECT  7.150 2.125 7.480 2.480 ;
        RECT  7.150 2.145 7.490 2.480 ;
        RECT  7.150 2.250 8.640 2.480 ;
        RECT  4.605 2.235 4.945 2.575 ;
        RECT  4.715 2.235 4.945 3.240 ;
        RECT  4.715 3.010 6.145 3.240 ;
        RECT  5.915 3.010 6.145 3.510 ;
        RECT  5.915 3.280 8.640 3.510 ;
        RECT  8.405 0.980 8.640 3.515 ;
        RECT  8.300 2.250 8.640 3.515 ;
        RECT  3.135 3.470 4.40 3.700 ;
        RECT  3.380 0.630 5.90 0.860 ;
        RECT  5.915 3.280 7.40 3.510 ;
    END
END DLLRQX2

MACRO DLLRQX1
    CLASS CORE ;
    FOREIGN DLLRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.480 1.615 3.035 2.060 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 2.970 1.240 3.780 ;
        RECT  0.900 0.700 1.240 1.040 ;
        RECT  0.900 0.700 1.135 3.780 ;
        RECT  0.755 2.250 1.135 2.630 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.840 2.095 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.500 7.530 1.840 ;
        RECT  7.055 1.500 7.435 2.635 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.945 -0.400 7.285 1.270 ;
        RECT  2.135 -0.400 2.475 0.710 ;
        RECT  0.180 -0.400 0.520 1.060 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.910 3.525 7.250 5.280 ;
        RECT  5.810 3.800 6.150 5.280 ;
        RECT  2.465 3.530 3.500 5.280 ;
        RECT  0.180 3.030 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.530 1.360 1.870 1.700 ;
        RECT  1.530 1.360 1.795 2.755 ;
        RECT  1.365 2.415 1.795 2.755 ;
        RECT  1.565 1.360 1.795 3.850 ;
        RECT  1.565 3.510 2.085 3.850 ;
        RECT  4.125 1.090 4.465 1.375 ;
        RECT  3.440 1.145 4.465 1.375 ;
        RECT  2.025 2.440 2.325 3.050 ;
        RECT  3.440 1.145 3.670 3.050 ;
        RECT  2.025 2.710 3.670 3.050 ;
        RECT  2.025 2.750 3.960 3.050 ;
        RECT  3.730 2.750 3.960 3.830 ;
        RECT  3.730 3.600 4.790 3.830 ;
        RECT  4.450 3.600 4.790 3.940 ;
        RECT  2.895 0.630 5.865 0.860 ;
        RECT  2.895 0.630 3.235 1.040 ;
        RECT  5.525 0.630 5.865 1.375 ;
        RECT  6.225 0.810 6.565 1.730 ;
        RECT  3.900 1.605 4.915 1.945 ;
        RECT  4.685 1.605 4.915 2.835 ;
        RECT  4.685 2.415 5.200 2.835 ;
        RECT  6.110 1.495 6.340 2.835 ;
        RECT  4.685 2.550 6.340 2.835 ;
        RECT  7.665 0.865 8.010 1.205 ;
        RECT  6.570 1.980 6.825 3.295 ;
        RECT  7.660 2.820 8.010 3.295 ;
        RECT  7.775 0.865 8.010 3.295 ;
        RECT  4.190 3.065 8.010 3.295 ;
        RECT  4.190 3.010 4.530 3.350 ;
        RECT  2.895 0.630 4.90 0.860 ;
        RECT  4.190 3.065 7.30 3.295 ;
    END
END DLLRQX1

MACRO DLLRQX0
    CLASS CORE ;
    FOREIGN DLLRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.640 2.110 2.110 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.350 0.660 1.160 1.000 ;
        RECT  0.125 2.800 0.795 3.240 ;
        RECT  0.350 0.660 0.580 3.240 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.345 3.240 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.230 6.245 2.755 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.310 -0.400 6.650 1.090 ;
        RECT  1.680 -0.400 2.020 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.410 3.965 6.590 5.280 ;
        RECT  1.955 3.660 3.195 5.280 ;
        RECT  0.455 3.600 0.795 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.810 1.360 1.150 2.570 ;
        RECT  2.440 2.200 2.725 2.570 ;
        RECT  0.810 2.340 2.725 2.570 ;
        RECT  1.025 2.340 1.255 4.000 ;
        RECT  1.025 3.660 1.495 4.000 ;
        RECT  2.955 1.200 3.850 1.540 ;
        RECT  2.955 1.200 3.185 3.240 ;
        RECT  2.385 2.860 3.185 3.240 ;
        RECT  1.485 3.010 3.770 3.240 ;
        RECT  1.485 3.010 1.775 3.420 ;
        RECT  3.540 3.010 3.770 4.250 ;
        RECT  3.540 3.965 4.395 4.250 ;
        RECT  2.480 0.630 5.250 0.970 ;
        RECT  4.910 0.630 5.250 1.540 ;
        RECT  5.610 0.630 5.950 2.000 ;
        RECT  5.610 1.770 6.865 2.000 ;
        RECT  6.560 1.770 6.865 2.365 ;
        RECT  6.560 1.770 6.790 3.275 ;
        RECT  5.650 2.985 6.790 3.275 ;
        RECT  7.070 1.360 7.380 1.665 ;
        RECT  3.415 1.770 3.700 2.540 ;
        RECT  4.460 2.200 4.800 2.540 ;
        RECT  3.415 2.310 4.800 2.540 ;
        RECT  4.075 2.310 4.305 3.735 ;
        RECT  7.040 3.140 7.380 3.735 ;
        RECT  7.095 1.360 7.380 3.735 ;
        RECT  4.075 3.505 7.380 3.735 ;
        RECT  1.485 3.010 2.20 3.240 ;
        RECT  2.480 0.630 4.80 0.970 ;
        RECT  4.075 3.505 6.60 3.735 ;
    END
END DLLRQX0

MACRO DLLQX4
    CLASS CORE ;
    FOREIGN DLLQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.645 1.550 1.135 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 1.130 8.695 3.880 ;
        RECT  6.860 2.180 8.695 2.410 ;
        RECT  6.860 1.130 7.200 3.880 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.470 ;
        RECT  6.100 -0.400 6.440 0.720 ;
        RECT  4.780 -0.400 5.120 0.985 ;
        RECT  2.460 -0.400 2.800 0.955 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 2.640 7.920 5.280 ;
        RECT  6.100 2.910 6.440 5.280 ;
        RECT  4.580 4.150 4.920 5.280 ;
        RECT  2.205 3.785 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  1.330 2.145 1.670 2.480 ;
        RECT  1.340 2.125 1.670 2.480 ;
        RECT  0.180 2.250 1.670 2.480 ;
        RECT  0.180 2.250 0.520 3.460 ;
        RECT  3.875 2.455 4.215 3.460 ;
        RECT  0.180 3.230 4.215 3.460 ;
        RECT  1.700 0.980 2.130 1.320 ;
        RECT  3.315 1.785 4.225 2.125 ;
        RECT  1.740 2.700 2.130 3.000 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.710 2.130 3.000 ;
        RECT  3.155 2.700 3.545 3.000 ;
        RECT  3.315 1.785 3.545 3.000 ;
        RECT  1.700 2.770 3.545 3.000 ;
        RECT  3.660 1.215 4.000 1.555 ;
        RECT  3.660 1.325 4.685 1.555 ;
        RECT  4.455 1.860 6.120 2.090 ;
        RECT  5.780 1.860 6.120 2.220 ;
        RECT  4.455 1.325 4.685 3.920 ;
        RECT  3.435 3.690 4.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  5.540 1.240 6.630 1.580 ;
        RECT  4.915 2.320 5.235 2.680 ;
        RECT  6.400 1.240 6.630 2.680 ;
        RECT  4.915 2.450 6.630 2.680 ;
        RECT  5.340 2.450 5.680 4.170 ;
        RECT  0.180 3.230 3.30 3.460 ;
    END
END DLLQX4

MACRO DLLQX2
    CLASS CORE ;
    FOREIGN DLLQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.615 5.160 2.080 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.550 6.915 2.020 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.240 1.140 3.480 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.320 ;
        RECT  4.900 -0.400 5.240 0.850 ;
        RECT  2.930 -0.400 3.270 0.810 ;
        RECT  0.240 -0.400 1.900 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.480 3.950 6.820 5.280 ;
        RECT  5.110 3.750 5.450 5.280 ;
        RECT  2.440 3.910 2.785 5.280 ;
        RECT  0.240 3.950 1.700 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.930 1.240 2.460 1.580 ;
        RECT  1.930 1.240 2.160 3.550 ;
        RECT  1.930 2.690 2.785 3.030 ;
        RECT  1.930 2.690 2.460 3.550 ;
        RECT  3.870 0.630 4.210 1.415 ;
        RECT  3.015 1.180 4.210 1.415 ;
        RECT  2.390 2.020 3.245 2.360 ;
        RECT  3.015 1.180 3.245 4.035 ;
        RECT  3.015 3.750 4.220 4.035 ;
        RECT  5.600 0.980 5.940 1.320 ;
        RECT  3.590 1.680 4.295 2.020 ;
        RECT  4.065 1.680 4.295 3.060 ;
        RECT  5.430 1.090 5.660 3.060 ;
        RECT  4.065 2.720 5.990 3.060 ;
        RECT  7.040 0.980 7.380 1.320 ;
        RECT  5.890 2.125 6.220 2.480 ;
        RECT  5.890 2.145 6.230 2.480 ;
        RECT  5.890 2.250 7.380 2.480 ;
        RECT  3.490 2.350 3.830 2.690 ;
        RECT  3.600 2.350 3.830 3.520 ;
        RECT  7.040 2.250 7.380 3.520 ;
        RECT  7.145 0.980 7.380 3.520 ;
        RECT  3.600 3.290 7.380 3.520 ;
        RECT  3.600 3.290 6.20 3.520 ;
    END
END DLLQX2

MACRO DLLQX1
    CLASS CORE ;
    FOREIGN DLLQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.945 2.970 1.285 3.780 ;
        RECT  0.945 0.700 1.285 1.040 ;
        RECT  0.945 0.700 1.175 3.780 ;
        RECT  0.755 2.250 1.175 2.630 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.210 2.095 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.500 6.900 1.840 ;
        RECT  6.425 1.500 6.805 2.125 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.315 -0.400 6.655 1.270 ;
        RECT  4.895 -0.400 5.235 1.375 ;
        RECT  1.795 -0.400 2.605 0.710 ;
        RECT  0.220 -0.400 0.565 1.040 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.280 3.525 6.620 5.280 ;
        RECT  5.180 3.800 5.520 5.280 ;
        RECT  2.465 3.530 2.870 5.280 ;
        RECT  0.220 2.970 0.565 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.515 1.360 1.870 1.700 ;
        RECT  1.515 1.360 1.795 3.850 ;
        RECT  1.515 2.940 1.805 3.850 ;
        RECT  1.515 3.510 2.085 3.850 ;
        RECT  3.495 1.035 3.835 1.375 ;
        RECT  2.810 1.145 3.835 1.375 ;
        RECT  2.810 1.145 3.040 2.545 ;
        RECT  2.025 2.205 3.040 2.545 ;
        RECT  2.025 2.245 3.330 2.545 ;
        RECT  3.100 2.245 3.330 3.830 ;
        RECT  3.100 3.600 4.160 3.830 ;
        RECT  3.820 3.600 4.160 3.940 ;
        RECT  5.595 0.810 5.935 1.150 ;
        RECT  3.270 1.605 4.285 1.945 ;
        RECT  4.055 1.605 4.285 2.835 ;
        RECT  4.055 2.415 4.570 2.835 ;
        RECT  5.480 0.905 5.710 2.835 ;
        RECT  4.055 2.550 5.710 2.835 ;
        RECT  7.035 0.865 7.380 1.205 ;
        RECT  5.940 1.980 6.195 3.295 ;
        RECT  7.030 2.820 7.380 3.295 ;
        RECT  7.145 0.865 7.380 3.295 ;
        RECT  3.560 3.065 7.380 3.295 ;
        RECT  3.560 3.010 3.900 3.350 ;
        RECT  3.560 3.065 6.50 3.295 ;
    END
END DLLQX1

MACRO DLLQX0
    CLASS CORE ;
    FOREIGN DLLQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.860 0.815 3.380 ;
        RECT  0.585 1.360 0.815 3.380 ;
        RECT  0.380 1.360 0.815 1.700 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.715 3.240 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.150 2.230 5.615 2.755 ;
        END
    END GN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.680 -0.400 6.020 1.090 ;
        RECT  4.280 -0.400 4.620 1.590 ;
        RECT  1.980 -0.400 2.320 0.980 ;
        RECT  0.380 -0.400 0.720 0.900 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.890 3.965 5.960 5.280 ;
        RECT  2.175 3.470 2.515 5.280 ;
        RECT  0.475 3.930 0.815 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.180 1.250 1.520 2.540 ;
        RECT  1.180 2.200 2.095 2.540 ;
        RECT  1.050 2.310 1.280 4.160 ;
        RECT  1.050 3.890 1.615 4.160 ;
        RECT  2.880 0.640 3.220 1.540 ;
        RECT  2.325 1.310 3.220 1.540 ;
        RECT  2.325 1.310 2.555 3.240 ;
        RECT  1.510 3.010 3.140 3.240 ;
        RECT  1.510 3.010 1.850 3.660 ;
        RECT  2.910 3.010 3.140 4.250 ;
        RECT  2.910 3.965 3.650 4.250 ;
        RECT  4.980 0.630 5.320 2.000 ;
        RECT  4.980 1.770 6.235 2.000 ;
        RECT  5.930 1.770 6.235 2.365 ;
        RECT  5.930 1.770 6.160 3.275 ;
        RECT  5.020 2.985 6.160 3.275 ;
        RECT  6.440 1.360 6.750 1.665 ;
        RECT  2.785 1.770 3.070 2.540 ;
        RECT  3.830 2.200 4.170 2.540 ;
        RECT  2.785 2.310 4.170 2.540 ;
        RECT  3.445 2.310 3.675 3.735 ;
        RECT  6.410 3.140 6.750 3.735 ;
        RECT  6.465 1.360 6.750 3.735 ;
        RECT  3.445 3.505 6.750 3.735 ;
        RECT  3.445 3.505 5.00 3.735 ;
    END
END DLLQX0

MACRO DLHX4
    CLASS CORE ;
    FOREIGN DLHX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.820 1.240 11.215 4.100 ;
        RECT  9.660 2.250 11.215 2.480 ;
        RECT  9.500 2.640 9.890 3.770 ;
        RECT  9.660 0.790 9.890 3.770 ;
        RECT  9.500 0.790 9.890 1.700 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.180 1.240 8.520 3.450 ;
        RECT  6.860 2.250 8.520 2.630 ;
        RECT  6.860 1.240 7.200 3.450 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.190 1.670 2.420 ;
        RECT  1.330 2.080 1.670 2.420 ;
        RECT  0.755 2.190 1.135 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.260 -0.400 10.600 0.720 ;
        RECT  6.100 -0.400 9.080 0.720 ;
        RECT  4.780 -0.400 5.120 0.995 ;
        RECT  2.460 -0.400 2.800 0.955 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  6.300 4.140 10.400 5.280 ;
        RECT  4.780 4.150 5.120 5.280 ;
        RECT  2.205 3.785 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  3.875 2.455 4.215 2.795 ;
        RECT  0.180 2.645 0.520 3.460 ;
        RECT  3.875 2.455 4.105 3.460 ;
        RECT  0.180 3.230 4.105 3.460 ;
        RECT  1.700 0.980 2.130 1.850 ;
        RECT  0.660 1.620 2.130 1.850 ;
        RECT  0.660 1.620 1.000 1.960 ;
        RECT  3.315 1.785 4.225 2.125 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.660 2.130 3.000 ;
        RECT  3.315 1.785 3.545 3.000 ;
        RECT  1.700 2.700 3.545 3.000 ;
        RECT  3.660 1.215 4.000 1.555 ;
        RECT  3.660 1.325 4.685 1.555 ;
        RECT  4.455 1.880 6.120 2.110 ;
        RECT  5.780 1.880 6.120 2.220 ;
        RECT  4.455 1.325 4.685 3.920 ;
        RECT  3.435 3.690 4.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  5.540 1.240 6.630 1.580 ;
        RECT  8.895 2.075 9.430 2.415 ;
        RECT  4.915 2.340 5.235 2.680 ;
        RECT  4.915 2.450 6.630 2.680 ;
        RECT  6.400 1.240 6.630 3.910 ;
        RECT  8.895 2.075 9.125 3.910 ;
        RECT  6.400 3.680 9.125 3.910 ;
        RECT  5.540 2.450 5.880 4.170 ;
        RECT  0.180 3.230 3.40 3.460 ;
        RECT  6.400 3.680 8.60 3.910 ;
    END
END DLHX4

MACRO DLHX2
    CLASS CORE ;
    FOREIGN DLHX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.240 1.135 3.480 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.785 1.615 6.445 2.080 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.240 2.400 3.480 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.190 8.065 2.635 ;
        RECT  7.150 2.190 8.065 2.420 ;
        RECT  7.150 2.080 7.490 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.320 ;
        RECT  6.160 -0.400 6.500 0.850 ;
        RECT  4.190 -0.400 4.530 0.810 ;
        RECT  0.180 -0.400 3.160 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.740 3.950 8.080 5.280 ;
        RECT  6.370 3.750 6.710 5.280 ;
        RECT  3.700 3.910 4.045 5.280 ;
        RECT  1.500 4.170 2.960 5.280 ;
        RECT  0.180 4.010 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.190 1.240 3.720 1.580 ;
        RECT  3.190 2.690 4.045 3.030 ;
        RECT  3.190 2.690 3.720 3.550 ;
        RECT  3.190 1.240 3.420 3.940 ;
        RECT  0.930 3.710 3.420 3.940 ;
        RECT  0.930 3.710 1.270 4.070 ;
        RECT  5.130 0.630 5.470 1.415 ;
        RECT  4.275 1.180 5.470 1.415 ;
        RECT  3.650 2.020 4.505 2.360 ;
        RECT  4.275 1.180 4.505 4.035 ;
        RECT  4.275 3.750 5.480 4.035 ;
        RECT  6.860 0.980 7.200 1.850 ;
        RECT  6.690 1.620 8.160 1.850 ;
        RECT  7.820 1.620 8.160 1.960 ;
        RECT  4.830 1.680 5.555 2.020 ;
        RECT  6.690 1.620 6.920 3.060 ;
        RECT  5.325 1.680 5.555 3.060 ;
        RECT  6.690 2.650 7.250 3.060 ;
        RECT  5.325 2.720 7.250 3.060 ;
        RECT  8.300 0.980 8.640 1.320 ;
        RECT  4.750 2.350 5.090 3.520 ;
        RECT  8.300 2.645 8.640 3.520 ;
        RECT  8.405 0.980 8.640 3.520 ;
        RECT  4.750 3.290 8.640 3.520 ;
        RECT  0.930 3.710 2.50 3.940 ;
        RECT  4.750 3.290 7.10 3.520 ;
    END
END DLHX2

MACRO DLHX1
    CLASS CORE ;
    FOREIGN DLHX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.820 0.520 3.880 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 2.970 1.960 3.780 ;
        RECT  1.535 0.700 1.960 1.040 ;
        RECT  1.535 0.700 1.765 3.215 ;
        RECT  1.385 2.250 1.765 2.630 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.840 2.095 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.075 7.435 2.635 ;
        RECT  6.570 2.075 7.435 2.320 ;
        RECT  6.570 1.980 6.855 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.945 -0.400 7.285 1.270 ;
        RECT  5.525 -0.400 5.865 1.375 ;
        RECT  2.425 -0.400 3.235 0.710 ;
        RECT  0.900 -0.400 1.240 1.060 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.910 3.525 7.250 5.280 ;
        RECT  5.810 3.800 6.150 5.280 ;
        RECT  3.095 3.530 3.500 5.280 ;
        RECT  0.900 3.030 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.160 1.360 2.500 1.700 ;
        RECT  2.160 1.360 2.425 2.350 ;
        RECT  1.995 2.010 2.425 2.350 ;
        RECT  2.195 1.360 2.425 3.850 ;
        RECT  2.195 3.510 2.715 3.850 ;
        RECT  3.440 1.035 4.465 1.375 ;
        RECT  3.440 1.035 3.670 2.780 ;
        RECT  2.655 2.440 3.670 2.780 ;
        RECT  2.655 2.480 3.960 2.780 ;
        RECT  3.730 2.480 3.960 3.940 ;
        RECT  3.730 3.600 4.790 3.940 ;
        RECT  6.225 0.810 6.565 1.730 ;
        RECT  6.110 1.500 7.530 1.730 ;
        RECT  7.190 1.500 7.530 1.840 ;
        RECT  3.900 1.605 4.915 1.945 ;
        RECT  4.685 1.605 4.915 2.835 ;
        RECT  4.685 2.415 5.200 2.835 ;
        RECT  6.110 1.495 6.340 2.835 ;
        RECT  4.685 2.550 6.435 2.835 ;
        RECT  7.665 0.865 8.010 1.205 ;
        RECT  7.660 2.820 8.010 3.295 ;
        RECT  7.775 0.865 8.010 3.295 ;
        RECT  4.190 3.065 8.010 3.295 ;
        RECT  4.190 3.010 4.530 3.350 ;
        RECT  4.190 3.065 7.40 3.295 ;
    END
END DLHX1

MACRO DLHX0
    CLASS CORE ;
    FOREIGN DLHX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.536  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.080 0.815 3.420 ;
        RECT  0.125 0.630 0.520 3.420 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.549  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.775 1.640 2.395 2.020 ;
        RECT  1.775 1.415 2.115 3.090 ;
        RECT  1.680 1.415 2.115 1.700 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.345 3.240 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.230 6.245 2.755 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.310 -0.400 6.650 1.090 ;
        RECT  4.910 -0.400 5.250 1.540 ;
        RECT  2.480 -0.400 2.820 0.970 ;
        RECT  0.880 -0.400 1.220 0.725 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.520 3.965 6.590 5.280 ;
        RECT  2.805 3.470 3.145 5.280 ;
        RECT  0.475 3.930 0.815 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.680 0.630 2.020 1.185 ;
        RECT  1.220 0.955 2.020 1.185 ;
        RECT  1.220 0.955 1.450 2.510 ;
        RECT  1.050 2.170 1.280 4.160 ;
        RECT  1.050 3.890 1.615 4.160 ;
        RECT  2.955 1.200 3.850 1.540 ;
        RECT  2.955 1.200 3.185 3.240 ;
        RECT  2.345 3.010 3.770 3.240 ;
        RECT  2.345 3.010 2.575 3.660 ;
        RECT  1.510 3.320 2.575 3.660 ;
        RECT  3.540 3.010 3.770 4.250 ;
        RECT  3.540 3.965 4.280 4.250 ;
        RECT  5.610 1.360 5.950 2.000 ;
        RECT  3.415 1.770 6.865 2.000 ;
        RECT  3.415 1.770 4.800 2.110 ;
        RECT  6.560 1.770 6.865 2.365 ;
        RECT  4.460 1.770 4.800 2.540 ;
        RECT  6.560 1.770 6.790 3.275 ;
        RECT  5.650 2.985 6.790 3.275 ;
        RECT  7.070 1.360 7.380 1.665 ;
        RECT  3.785 2.440 4.230 2.780 ;
        RECT  4.000 2.440 4.230 3.735 ;
        RECT  7.040 3.095 7.380 3.735 ;
        RECT  7.095 1.360 7.380 3.735 ;
        RECT  4.000 3.505 7.380 3.735 ;
        RECT  3.415 1.770 5.60 2.000 ;
        RECT  4.000 3.505 6.40 3.735 ;
    END
END DLHX0

MACRO DLHSX4
    CLASS CORE ;
    FOREIGN DLHSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.070 1.240 10.410 3.450 ;
        RECT  8.750 2.250 10.410 2.630 ;
        RECT  8.750 1.240 9.090 3.450 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.805 1.640 4.285 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 1.240 13.105 4.100 ;
        RECT  11.550 2.250 13.105 2.480 ;
        RECT  11.390 2.640 11.780 3.770 ;
        RECT  11.550 0.790 11.780 3.770 ;
        RECT  11.390 0.790 11.780 1.700 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.980 2.250 5.545 2.635 ;
        RECT  4.980 2.080 5.310 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  12.150 -0.400 12.490 0.720 ;
        RECT  6.870 -0.400 10.970 0.720 ;
        RECT  5.450 -0.400 5.790 1.320 ;
        RECT  4.030 -0.400 4.370 0.970 ;
        RECT  1.770 -0.400 2.110 0.950 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  7.990 4.140 12.290 5.280 ;
        RECT  6.740 2.640 7.050 5.280 ;
        RECT  5.170 3.625 5.510 5.280 ;
        RECT  3.925 3.900 4.265 5.280 ;
        RECT  1.540 4.110 1.880 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.765 1.410 ;
        RECT  1.535 1.180 1.765 2.090 ;
        RECT  1.535 1.805 1.875 2.090 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  2.110 1.235 3.140 1.575 ;
        RECT  2.110 1.235 2.340 2.550 ;
        RECT  1.845 2.320 2.340 2.550 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.845 2.320 2.075 3.610 ;
        RECT  0.170 3.380 2.340 3.610 ;
        RECT  2.110 3.380 2.340 3.965 ;
        RECT  2.110 3.625 3.035 3.965 ;
        RECT  4.730 0.980 5.070 1.850 ;
        RECT  4.520 1.620 6.030 1.850 ;
        RECT  5.690 1.620 6.030 1.960 ;
        RECT  4.520 1.620 4.750 2.935 ;
        RECT  3.030 2.595 4.750 2.935 ;
        RECT  6.170 0.980 6.510 1.320 ;
        RECT  3.235 1.805 3.575 2.145 ;
        RECT  2.570 1.915 3.575 2.145 ;
        RECT  6.275 0.980 6.510 2.420 ;
        RECT  5.930 2.190 6.510 2.420 ;
        RECT  2.305 2.780 2.800 3.080 ;
        RECT  2.570 1.915 2.800 3.395 ;
        RECT  2.570 3.165 6.270 3.395 ;
        RECT  5.930 2.190 6.270 3.550 ;
        RECT  10.785 2.075 11.320 2.415 ;
        RECT  7.430 1.240 7.770 3.910 ;
        RECT  10.785 2.075 11.015 3.910 ;
        RECT  7.430 3.680 11.015 3.910 ;
        RECT  0.170 3.380 1.80 3.610 ;
        RECT  2.570 3.165 5.40 3.395 ;
        RECT  7.430 3.680 10.40 3.910 ;
    END
END DLHSX4

MACRO DLHSX2
    CLASS CORE ;
    FOREIGN DLHSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 1.240 8.065 3.480 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.795 2.130 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 1.640 1.135 2.465 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 1.240 9.340 3.480 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.190 5.545 2.635 ;
        RECT  4.505 2.190 5.545 2.420 ;
        RECT  4.505 2.080 4.845 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  6.920 -0.400 9.900 0.720 ;
        RECT  4.940 -0.400 5.280 1.320 ;
        RECT  3.445 -0.400 3.785 0.955 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.560 4.010 9.900 5.280 ;
        RECT  7.120 4.170 8.580 5.280 ;
        RECT  5.025 3.700 5.365 5.280 ;
        RECT  3.850 3.875 4.190 5.280 ;
        RECT  1.440 4.170 1.780 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.950 ;
        RECT  0.180 0.630 0.410 2.925 ;
        RECT  1.365 1.890 1.650 2.925 ;
        RECT  0.180 2.695 1.650 2.925 ;
        RECT  0.740 2.695 1.080 3.150 ;
        RECT  2.245 1.270 2.585 1.610 ;
        RECT  1.880 1.380 2.585 1.610 ;
        RECT  0.170 3.155 0.510 3.610 ;
        RECT  0.170 3.380 2.110 3.610 ;
        RECT  1.880 1.380 2.110 3.935 ;
        RECT  1.880 3.705 2.960 3.935 ;
        RECT  2.620 3.705 2.960 4.240 ;
        RECT  1.965 0.680 2.305 1.040 ;
        RECT  1.965 0.810 3.045 1.040 ;
        RECT  4.220 0.980 4.560 1.850 ;
        RECT  4.025 1.620 5.645 1.850 ;
        RECT  5.305 1.620 5.645 1.960 ;
        RECT  4.025 1.620 4.255 3.010 ;
        RECT  2.815 0.810 3.045 3.010 ;
        RECT  2.815 2.670 3.240 3.010 ;
        RECT  4.025 2.650 4.605 3.010 ;
        RECT  2.815 2.780 4.605 3.010 ;
        RECT  5.660 0.980 6.125 1.320 ;
        RECT  2.340 2.090 2.585 3.470 ;
        RECT  5.785 2.645 6.125 3.470 ;
        RECT  5.890 0.980 6.125 3.470 ;
        RECT  2.340 3.240 6.125 3.470 ;
        RECT  6.360 1.170 6.700 3.940 ;
        RECT  6.360 3.710 9.150 3.940 ;
        RECT  8.810 3.710 9.150 4.070 ;
        RECT  2.340 3.240 5.30 3.470 ;
        RECT  6.360 3.710 8.20 3.940 ;
    END
END DLHSX2

MACRO DLHSX1
    CLASS CORE ;
    FOREIGN DLHSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.235 2.250 8.695 2.630 ;
        RECT  8.235 0.700 8.465 3.515 ;
        RECT  8.120 3.270 8.460 4.080 ;
        RECT  8.120 0.700 8.465 1.040 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.560 0.820 9.955 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.655 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.142  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.860 2.030 3.260 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.075 6.175 2.635 ;
        RECT  5.345 2.075 6.175 2.320 ;
        RECT  5.345 1.760 5.630 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.840 -0.400 9.180 1.060 ;
        RECT  7.320 -0.400 7.660 0.710 ;
        RECT  5.665 -0.400 6.005 0.665 ;
        RECT  4.165 -0.400 4.505 1.340 ;
        RECT  1.480 -0.400 1.820 1.180 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.840 3.330 9.180 5.280 ;
        RECT  7.185 4.170 7.525 5.280 ;
        RECT  5.885 3.525 6.225 5.280 ;
        RECT  4.570 3.525 4.910 5.280 ;
        RECT  1.750 3.840 2.095 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 1.210 0.520 1.895 ;
        RECT  0.170 1.555 2.155 1.895 ;
        RECT  0.170 1.210 0.400 3.250 ;
        RECT  0.170 3.020 1.120 3.250 ;
        RECT  0.890 3.020 1.120 4.175 ;
        RECT  0.890 3.835 1.280 4.175 ;
        RECT  2.430 1.250 3.105 1.590 ;
        RECT  0.630 2.155 2.660 2.495 ;
        RECT  2.430 1.250 2.660 3.845 ;
        RECT  2.430 3.525 3.510 3.845 ;
        RECT  4.885 0.810 5.245 1.150 ;
        RECT  2.485 0.630 3.675 0.970 ;
        RECT  4.885 0.895 6.325 1.150 ;
        RECT  6.035 0.895 6.325 1.840 ;
        RECT  6.035 1.500 6.375 1.840 ;
        RECT  3.445 0.630 3.675 2.835 ;
        RECT  4.885 0.810 5.115 2.835 ;
        RECT  3.445 2.470 5.115 2.835 ;
        RECT  3.445 2.550 5.410 2.835 ;
        RECT  6.600 0.980 6.985 1.320 ;
        RECT  2.890 2.680 3.215 3.295 ;
        RECT  6.635 2.720 6.985 3.295 ;
        RECT  6.750 0.980 6.985 3.295 ;
        RECT  2.890 3.065 6.985 3.295 ;
        RECT  7.300 1.170 7.750 1.510 ;
        RECT  7.300 2.130 7.985 2.505 ;
        RECT  7.300 1.170 7.530 3.820 ;
        RECT  7.185 3.445 7.530 3.820 ;
        RECT  0.630 2.155 1.80 2.495 ;
        RECT  2.890 3.065 5.80 3.295 ;
    END
END DLHSX1

MACRO DLHSX0
    CLASS CORE ;
    FOREIGN DLHSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.481  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.595 2.250 7.435 2.630 ;
        RECT  6.595 0.675 7.240 1.015 ;
        RECT  6.180 3.965 6.825 4.250 ;
        RECT  6.595 0.675 6.825 4.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.559  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 0.630 8.705 4.135 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.460 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.760 1.765 3.350 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.930 2.230 5.270 2.755 ;
        RECT  4.535 2.230 5.270 2.630 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.595 -0.400 7.940 0.970 ;
        RECT  5.450 -0.400 6.365 1.145 ;
        RECT  3.950 -0.400 4.290 1.540 ;
        RECT  1.320 -0.400 1.660 1.460 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.055 3.885 7.865 5.280 ;
        RECT  4.560 3.965 5.630 5.280 ;
        RECT  1.755 3.580 2.095 5.280 ;
        RECT  0.180 3.930 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.990 ;
        RECT  0.115 1.760 1.765 1.990 ;
        RECT  1.425 1.760 1.765 2.070 ;
        RECT  0.115 0.630 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  1.995 1.230 2.890 1.540 ;
        RECT  0.575 2.300 2.225 2.530 ;
        RECT  0.575 2.300 0.915 2.955 ;
        RECT  1.995 1.230 2.225 3.240 ;
        RECT  1.995 3.010 2.810 3.240 ;
        RECT  2.580 3.010 2.810 4.250 ;
        RECT  2.580 3.965 3.320 4.250 ;
        RECT  4.650 1.385 4.990 2.000 ;
        RECT  2.455 1.770 5.905 2.000 ;
        RECT  2.455 1.770 2.740 2.110 ;
        RECT  5.600 1.770 5.905 2.365 ;
        RECT  3.500 1.770 3.840 2.635 ;
        RECT  3.500 1.770 3.800 2.655 ;
        RECT  5.600 1.770 5.830 3.275 ;
        RECT  4.690 2.985 5.830 3.275 ;
        RECT  2.825 2.440 3.270 2.780 ;
        RECT  3.040 2.440 3.270 3.735 ;
        RECT  6.080 3.095 6.365 3.735 ;
        RECT  6.135 1.505 6.365 3.735 ;
        RECT  3.040 3.505 6.365 3.735 ;
        RECT  7.055 1.375 7.895 1.715 ;
        RECT  7.665 2.395 8.070 2.735 ;
        RECT  7.665 1.375 7.895 3.335 ;
        RECT  7.155 2.995 7.895 3.335 ;
        RECT  2.455 1.770 4.80 2.000 ;
        RECT  3.040 3.505 5.30 3.735 ;
    END
END DLHSX0

MACRO DLHSQX4
    CLASS CORE ;
    FOREIGN DLHSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.805 1.640 4.285 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.200 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 1.130 10.585 3.880 ;
        RECT  8.910 2.130 10.585 2.360 ;
        RECT  8.750 2.640 9.140 3.880 ;
        RECT  8.910 1.130 9.140 3.880 ;
        RECT  8.750 1.130 9.140 1.470 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.980 2.250 5.545 2.635 ;
        RECT  4.980 2.080 5.310 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.470 ;
        RECT  6.870 -0.400 8.330 0.720 ;
        RECT  5.450 -0.400 5.790 1.320 ;
        RECT  4.030 -0.400 4.370 0.970 ;
        RECT  1.770 -0.400 2.110 0.950 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 2.640 9.810 5.280 ;
        RECT  7.990 3.950 8.330 5.280 ;
        RECT  6.740 2.640 7.050 5.280 ;
        RECT  5.170 3.625 5.510 5.280 ;
        RECT  3.925 3.900 4.265 5.280 ;
        RECT  1.540 4.110 1.880 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.875 1.410 ;
        RECT  1.535 1.180 1.875 2.090 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  2.110 1.235 3.140 1.575 ;
        RECT  2.110 1.235 2.340 2.550 ;
        RECT  1.845 2.320 2.340 2.550 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.845 2.320 2.075 3.610 ;
        RECT  0.170 3.380 2.340 3.610 ;
        RECT  2.110 3.380 2.340 3.855 ;
        RECT  2.110 3.625 3.035 3.855 ;
        RECT  2.695 3.625 3.035 3.965 ;
        RECT  4.730 0.980 5.070 1.850 ;
        RECT  4.520 1.620 6.030 1.850 ;
        RECT  5.690 1.620 6.030 1.960 ;
        RECT  4.520 1.620 4.750 2.935 ;
        RECT  3.030 2.595 4.750 2.935 ;
        RECT  6.170 0.980 6.510 1.320 ;
        RECT  3.235 1.805 3.575 2.145 ;
        RECT  2.570 1.915 3.575 2.145 ;
        RECT  2.305 2.780 2.800 3.080 ;
        RECT  2.570 1.915 2.800 3.395 ;
        RECT  2.570 3.165 6.510 3.395 ;
        RECT  6.275 0.980 6.510 3.550 ;
        RECT  5.930 2.645 6.510 3.550 ;
        RECT  7.430 2.075 8.680 2.415 ;
        RECT  7.430 1.240 7.770 3.550 ;
        RECT  0.170 3.380 1.70 3.610 ;
        RECT  2.570 3.165 5.30 3.395 ;
    END
END DLHSQX4

MACRO DLHSQX2
    CLASS CORE ;
    FOREIGN DLHSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.680 2.640 8.070 3.480 ;
        RECT  7.840 1.240 8.070 3.480 ;
        RECT  7.680 1.240 8.070 1.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.795 2.130 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.690 1.640 1.135 2.465 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.190 5.545 2.635 ;
        RECT  4.505 2.190 5.545 2.420 ;
        RECT  4.505 2.080 4.845 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.920 -0.400 8.580 0.720 ;
        RECT  4.940 -0.400 5.280 1.320 ;
        RECT  3.445 -0.400 3.785 0.955 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.120 4.170 8.580 5.280 ;
        RECT  5.025 3.700 5.365 5.280 ;
        RECT  3.850 3.875 4.190 5.280 ;
        RECT  1.440 4.170 1.780 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.950 ;
        RECT  0.180 0.630 0.410 2.925 ;
        RECT  1.365 1.890 1.650 2.925 ;
        RECT  0.180 2.695 1.650 2.925 ;
        RECT  0.740 2.695 1.080 3.150 ;
        RECT  1.880 1.270 2.585 1.610 ;
        RECT  0.170 3.155 0.510 3.610 ;
        RECT  0.170 3.380 2.110 3.610 ;
        RECT  1.880 1.270 2.110 3.935 ;
        RECT  1.880 3.705 2.960 3.935 ;
        RECT  2.620 3.705 2.960 4.240 ;
        RECT  1.965 0.680 3.045 1.020 ;
        RECT  4.220 0.980 4.560 1.850 ;
        RECT  4.025 1.620 5.645 1.850 ;
        RECT  5.305 1.620 5.645 1.960 ;
        RECT  4.025 1.620 4.255 3.010 ;
        RECT  2.815 0.680 3.045 3.010 ;
        RECT  4.025 2.650 4.605 3.010 ;
        RECT  2.815 2.670 4.605 3.010 ;
        RECT  5.660 0.980 6.125 1.320 ;
        RECT  2.340 2.090 2.585 3.470 ;
        RECT  5.785 2.645 6.125 3.470 ;
        RECT  5.890 0.980 6.125 3.470 ;
        RECT  2.340 3.240 6.125 3.470 ;
        RECT  6.360 1.880 7.610 2.220 ;
        RECT  6.360 1.170 6.700 3.540 ;
        RECT  2.340 3.240 5.70 3.470 ;
    END
END DLHSQX2

MACRO DLHSQX1
    CLASS CORE ;
    FOREIGN DLHSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 3.270 8.695 4.180 ;
        RECT  8.465 0.820 8.695 4.180 ;
        RECT  8.300 0.820 8.695 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.510 4.350 2.220 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.142  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.860 1.975 3.270 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.980 5.545 2.635 ;
        RECT  5.055 1.980 5.545 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.060 ;
        RECT  5.330 -0.400 5.670 1.175 ;
        RECT  3.870 -0.400 4.210 1.280 ;
        RECT  1.210 -0.400 1.550 0.715 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 3.330 7.920 5.280 ;
        RECT  5.400 3.525 5.740 5.280 ;
        RECT  4.290 3.825 4.630 5.280 ;
        RECT  1.655 3.840 1.975 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.120 1.035 0.520 1.465 ;
        RECT  0.120 1.235 1.970 1.465 ;
        RECT  1.630 1.235 1.970 2.170 ;
        RECT  0.120 1.035 0.350 3.250 ;
        RECT  0.120 3.020 1.120 3.250 ;
        RECT  0.890 3.020 1.120 4.175 ;
        RECT  0.890 3.835 1.280 4.175 ;
        RECT  2.205 1.250 2.810 1.590 ;
        RECT  0.580 2.290 0.865 2.630 ;
        RECT  0.580 2.400 2.435 2.630 ;
        RECT  2.205 1.250 2.435 4.115 ;
        RECT  2.205 3.775 3.230 4.115 ;
        RECT  2.190 0.630 3.530 0.970 ;
        RECT  4.580 0.810 4.950 1.730 ;
        RECT  4.580 1.500 6.035 1.730 ;
        RECT  5.740 1.500 6.035 1.840 ;
        RECT  3.300 0.630 3.530 2.835 ;
        RECT  3.300 2.470 3.640 2.835 ;
        RECT  4.580 0.810 4.810 2.835 ;
        RECT  3.300 2.550 4.925 2.835 ;
        RECT  6.045 0.900 6.500 1.240 ;
        RECT  2.665 2.950 2.950 3.295 ;
        RECT  6.150 2.540 6.500 3.295 ;
        RECT  2.665 3.065 6.500 3.295 ;
        RECT  6.265 0.900 6.500 3.350 ;
        RECT  6.160 2.540 6.500 3.350 ;
        RECT  6.780 0.940 7.155 4.180 ;
        RECT  6.780 2.160 8.160 2.500 ;
        RECT  6.780 2.160 7.160 4.180 ;
        RECT  2.665 3.065 5.10 3.295 ;
    END
END DLHSQX1

MACRO DLHSQX0
    CLASS CORE ;
    FOREIGN DLHSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.555 2.995 8.075 3.335 ;
        RECT  7.845 1.260 8.075 3.335 ;
        RECT  7.665 1.260 8.075 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.460 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.760 1.765 3.350 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.930 2.230 5.270 2.755 ;
        RECT  4.535 2.230 5.270 2.630 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.595 -0.400 7.940 0.900 ;
        RECT  5.450 -0.400 6.365 1.145 ;
        RECT  3.950 -0.400 4.290 1.540 ;
        RECT  1.320 -0.400 1.660 1.460 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.055 3.795 7.840 5.280 ;
        RECT  4.450 3.965 5.630 5.280 ;
        RECT  1.755 3.580 2.095 5.280 ;
        RECT  0.180 3.930 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.990 ;
        RECT  0.115 1.760 1.765 1.990 ;
        RECT  1.425 1.760 1.765 2.070 ;
        RECT  0.115 0.630 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  1.995 1.230 2.890 1.540 ;
        RECT  0.575 2.300 2.225 2.530 ;
        RECT  0.575 2.300 0.915 2.955 ;
        RECT  1.995 1.230 2.225 3.240 ;
        RECT  1.995 3.010 2.810 3.240 ;
        RECT  2.580 3.010 2.810 4.250 ;
        RECT  2.580 3.965 3.320 4.250 ;
        RECT  4.650 1.385 4.990 2.000 ;
        RECT  2.455 1.770 5.905 2.000 ;
        RECT  2.455 1.770 2.740 2.110 ;
        RECT  5.600 1.770 5.905 2.365 ;
        RECT  3.500 1.770 3.840 2.635 ;
        RECT  3.500 1.770 3.800 2.655 ;
        RECT  5.600 1.770 5.830 3.275 ;
        RECT  4.690 2.985 5.830 3.275 ;
        RECT  2.825 2.440 3.270 2.780 ;
        RECT  3.040 2.440 3.270 3.735 ;
        RECT  6.080 3.095 6.365 3.735 ;
        RECT  6.135 1.505 6.365 3.735 ;
        RECT  3.040 3.505 6.365 3.735 ;
        RECT  6.595 0.655 7.220 0.995 ;
        RECT  6.595 2.275 7.615 2.615 ;
        RECT  6.595 0.655 6.825 4.250 ;
        RECT  6.180 3.965 6.825 4.250 ;
        RECT  2.455 1.770 4.30 2.000 ;
        RECT  3.040 3.505 5.20 3.735 ;
    END
END DLHSQX0

MACRO DLHRX4
    CLASS CORE ;
    FOREIGN DLHRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 1.240 13.105 4.100 ;
        RECT  11.550 2.250 13.105 2.480 ;
        RECT  11.390 2.640 11.780 3.770 ;
        RECT  11.550 0.790 11.780 3.770 ;
        RECT  11.390 0.790 11.780 1.700 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.900 3.025 6.280 3.385 ;
        RECT  5.780 2.855 6.240 3.260 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.070 1.240 10.410 3.450 ;
        RECT  8.750 2.250 10.410 2.630 ;
        RECT  8.750 1.240 9.090 3.450 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.190 1.670 2.420 ;
        RECT  1.330 2.080 1.670 2.420 ;
        RECT  0.755 2.190 1.135 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  12.150 -0.400 12.490 0.720 ;
        RECT  6.870 -0.400 10.970 0.720 ;
        RECT  5.450 -0.400 5.790 1.205 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  7.990 4.140 12.290 5.280 ;
        RECT  6.670 2.925 7.010 5.280 ;
        RECT  4.545 4.150 4.885 5.280 ;
        RECT  2.205 3.900 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  0.180 2.645 0.520 3.460 ;
        RECT  3.875 2.455 4.215 3.460 ;
        RECT  0.180 3.230 4.215 3.460 ;
        RECT  1.700 0.980 2.130 1.850 ;
        RECT  0.660 1.620 2.130 1.850 ;
        RECT  0.660 1.620 1.000 1.960 ;
        RECT  3.315 1.785 4.225 2.125 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.660 2.130 3.000 ;
        RECT  3.315 1.785 3.545 3.000 ;
        RECT  1.700 2.700 3.545 3.000 ;
        RECT  2.460 0.630 5.145 0.955 ;
        RECT  4.915 0.630 5.145 1.665 ;
        RECT  6.170 0.950 6.510 1.665 ;
        RECT  4.915 1.435 6.510 1.665 ;
        RECT  3.660 1.215 4.685 1.555 ;
        RECT  4.455 1.895 7.200 2.125 ;
        RECT  6.860 1.895 7.200 2.235 ;
        RECT  4.455 1.215 4.685 3.920 ;
        RECT  4.455 3.580 5.685 3.920 ;
        RECT  3.435 3.690 5.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  10.785 2.075 11.320 2.415 ;
        RECT  4.915 2.355 6.630 2.585 ;
        RECT  4.915 2.355 5.200 2.695 ;
        RECT  6.410 2.465 7.770 2.695 ;
        RECT  7.430 1.240 7.770 3.910 ;
        RECT  10.785 2.075 11.015 3.910 ;
        RECT  7.430 3.680 11.015 3.910 ;
        RECT  0.180 3.230 3.80 3.460 ;
        RECT  2.460 0.630 4.60 0.955 ;
        RECT  4.455 1.895 6.60 2.125 ;
        RECT  3.435 3.690 4.90 3.920 ;
        RECT  7.430 3.680 10.80 3.910 ;
    END
END DLHRX4

MACRO DLHRX2
    CLASS CORE ;
    FOREIGN DLHRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.240 1.135 3.480 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.400 2.595 4.915 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.015 1.640 7.575 2.085 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.240 2.400 3.480 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.190 9.325 2.635 ;
        RECT  8.410 2.190 9.325 2.420 ;
        RECT  8.410 2.080 8.750 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.800 -0.400 9.140 1.320 ;
        RECT  0.180 -0.400 4.220 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.800 3.680 9.140 5.280 ;
        RECT  7.485 3.680 7.825 5.280 ;
        RECT  5.195 3.930 5.535 5.280 ;
        RECT  1.500 4.170 2.960 5.280 ;
        RECT  0.180 4.010 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  3.270 1.240 3.720 1.795 ;
        RECT  3.270 1.565 5.115 1.795 ;
        RECT  4.830 1.565 5.115 1.905 ;
        RECT  3.270 2.640 3.720 3.550 ;
        RECT  3.270 1.240 3.500 3.940 ;
        RECT  0.930 3.710 3.500 3.940 ;
        RECT  0.930 3.710 1.270 4.070 ;
        RECT  5.345 1.090 6.210 1.335 ;
        RECT  3.730 2.025 4.070 2.365 ;
        RECT  3.730 2.135 5.575 2.365 ;
        RECT  5.345 1.090 5.575 3.700 ;
        RECT  4.395 3.470 6.595 3.700 ;
        RECT  4.395 3.470 4.735 3.810 ;
        RECT  6.255 3.470 6.595 3.810 ;
        RECT  4.640 0.630 7.530 0.860 ;
        RECT  7.300 0.630 7.530 1.310 ;
        RECT  4.640 0.630 4.980 1.215 ;
        RECT  7.300 0.970 7.640 1.310 ;
        RECT  7.950 0.980 8.380 1.850 ;
        RECT  7.950 1.620 9.420 1.850 ;
        RECT  5.805 1.565 6.765 1.905 ;
        RECT  9.080 1.620 9.420 1.960 ;
        RECT  6.535 1.565 6.765 2.780 ;
        RECT  7.950 0.980 8.180 2.990 ;
        RECT  6.535 2.480 8.180 2.780 ;
        RECT  7.950 2.650 8.380 2.990 ;
        RECT  9.560 0.980 9.900 1.320 ;
        RECT  5.865 2.235 6.205 2.575 ;
        RECT  5.975 2.235 6.205 3.240 ;
        RECT  5.975 3.010 7.405 3.240 ;
        RECT  7.175 3.220 9.900 3.450 ;
        RECT  9.665 0.980 9.900 3.455 ;
        RECT  9.560 2.645 9.900 3.455 ;
        RECT  0.930 3.710 2.20 3.940 ;
        RECT  4.395 3.470 5.80 3.700 ;
        RECT  4.640 0.630 6.30 0.860 ;
        RECT  7.175 3.220 8.70 3.450 ;
    END
END DLHRX2

MACRO DLHRX1
    CLASS CORE ;
    FOREIGN DLHRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.620 2.970 1.960 3.780 ;
        RECT  1.470 0.700 1.960 1.040 ;
        RECT  1.470 0.700 1.765 3.215 ;
        RECT  1.385 2.250 1.765 2.630 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.110 1.615 3.665 2.060 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.820 0.520 3.880 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.470 2.095 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.075 8.065 2.635 ;
        RECT  7.200 2.075 8.065 2.320 ;
        RECT  7.200 1.980 7.485 2.320 ;
        END
    END G
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.540 3.525 7.880 5.280 ;
        RECT  6.440 3.800 6.780 5.280 ;
        RECT  3.095 3.530 4.130 5.280 ;
        RECT  0.900 3.030 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.575 -0.400 7.915 1.270 ;
        RECT  2.765 -0.400 3.105 0.710 ;
        RECT  0.900 -0.400 1.240 1.060 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.160 1.360 2.500 1.700 ;
        RECT  2.160 1.360 2.425 2.350 ;
        RECT  1.995 2.010 2.425 2.350 ;
        RECT  2.195 1.360 2.425 3.850 ;
        RECT  2.195 3.510 2.715 3.850 ;
        RECT  4.755 1.090 5.095 1.375 ;
        RECT  4.070 1.145 5.095 1.375 ;
        RECT  2.655 2.440 2.955 3.050 ;
        RECT  4.070 1.145 4.300 3.050 ;
        RECT  2.655 2.710 4.300 3.050 ;
        RECT  2.655 2.750 4.590 3.050 ;
        RECT  4.360 2.750 4.590 3.940 ;
        RECT  4.360 3.600 5.420 3.940 ;
        RECT  3.525 0.630 6.495 0.860 ;
        RECT  3.525 0.630 3.865 1.040 ;
        RECT  6.155 0.630 6.495 1.375 ;
        RECT  6.855 0.810 7.195 1.730 ;
        RECT  6.740 1.500 8.160 1.730 ;
        RECT  7.820 1.500 8.160 1.840 ;
        RECT  4.530 1.605 5.545 1.945 ;
        RECT  5.315 1.605 5.545 2.835 ;
        RECT  5.315 2.415 5.830 2.835 ;
        RECT  6.740 1.495 6.970 2.835 ;
        RECT  5.315 2.550 7.065 2.835 ;
        RECT  8.295 0.865 8.640 1.205 ;
        RECT  8.290 2.820 8.640 3.295 ;
        RECT  8.405 0.865 8.640 3.295 ;
        RECT  4.820 3.065 8.640 3.295 ;
        RECT  4.820 3.010 5.160 3.350 ;
        RECT  3.525 0.630 5.30 0.860 ;
        RECT  4.820 3.065 7.70 3.295 ;
    END
END DLHRX1

MACRO DLHRX0
    CLASS CORE ;
    FOREIGN DLHRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.910 1.890 5.545 2.630 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.469  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.925 3.130 7.445 3.470 ;
        RECT  7.215 0.630 7.445 3.470 ;
        RECT  7.055 2.250 7.445 2.630 ;
        RECT  6.690 0.630 7.445 0.960 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.443  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.880 6.175 3.170 ;
        RECT  5.775 1.030 6.175 1.410 ;
        RECT  5.775 1.030 6.005 3.170 ;
        RECT  5.260 1.250 6.005 1.605 ;
        END
    END QN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.180 2.595 2.630 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 2.190 1.765 2.630 ;
        END
    END G
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.925 3.930 7.265 5.280 ;
        RECT  4.110 3.860 5.330 5.280 ;
        RECT  0.880 3.565 1.820 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.210 -0.400 6.205 0.800 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.720 0.520 1.170 ;
        RECT  1.610 0.630 1.950 1.170 ;
        RECT  0.115 0.940 1.950 1.170 ;
        RECT  0.115 0.720 0.345 4.055 ;
        RECT  0.115 3.715 0.520 4.055 ;
        RECT  0.750 1.400 1.820 1.700 ;
        RECT  0.575 1.935 0.980 2.275 ;
        RECT  0.750 1.400 0.980 3.090 ;
        RECT  3.625 1.805 3.965 3.090 ;
        RECT  0.750 2.860 3.965 3.090 ;
        RECT  2.430 2.860 2.770 3.190 ;
        RECT  1.480 2.860 1.820 3.205 ;
        RECT  2.180 0.680 4.750 0.910 ;
        RECT  2.180 0.680 2.520 1.020 ;
        RECT  4.410 0.680 4.750 1.035 ;
        RECT  3.380 1.195 3.720 1.535 ;
        RECT  3.380 1.305 4.540 1.535 ;
        RECT  4.310 1.305 4.540 3.630 ;
        RECT  4.310 2.985 4.730 3.630 ;
        RECT  2.880 3.400 6.235 3.630 ;
        RECT  5.910 3.400 6.235 3.750 ;
        RECT  2.880 3.400 3.220 3.885 ;
        RECT  6.465 1.320 6.985 1.660 ;
        RECT  6.235 2.305 6.695 2.645 ;
        RECT  6.465 1.320 6.695 4.250 ;
        RECT  6.035 3.980 6.695 4.250 ;
        RECT  0.750 2.860 2.90 3.090 ;
        RECT  2.180 0.680 3.70 0.910 ;
        RECT  2.880 3.400 5.80 3.630 ;
    END
END DLHRX0

MACRO DLHRSX4
    CLASS CORE ;
    FOREIGN DLHRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.782  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.330 1.240 11.670 3.450 ;
        RECT  10.010 2.250 11.670 2.630 ;
        RECT  10.010 1.240 10.350 3.450 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.140 2.030 2.480 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.140 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.065 1.640 5.545 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 1.240 14.365 4.100 ;
        RECT  12.810 2.250 14.365 2.480 ;
        RECT  12.650 2.640 13.040 3.770 ;
        RECT  12.810 0.790 13.040 3.770 ;
        RECT  12.650 0.790 13.040 1.700 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.240 2.250 6.805 2.635 ;
        RECT  6.240 2.080 6.570 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.410 -0.400 13.750 0.720 ;
        RECT  8.130 -0.400 12.230 0.720 ;
        RECT  6.710 -0.400 7.050 1.320 ;
        RECT  2.330 -0.400 2.670 0.655 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  9.250 4.140 13.550 5.280 ;
        RECT  8.000 2.640 8.310 5.280 ;
        RECT  6.430 3.625 6.770 5.280 ;
        RECT  5.185 3.900 5.525 5.280 ;
        RECT  1.540 3.930 2.920 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.910 ;
        RECT  1.365 1.680 2.730 1.910 ;
        RECT  2.500 1.680 2.730 2.610 ;
        RECT  2.510 2.290 2.840 2.625 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  4.060 1.235 4.400 1.575 ;
        RECT  3.070 1.345 4.400 1.575 ;
        RECT  1.995 2.740 2.310 3.700 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.995 2.775 2.335 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 3.525 3.700 ;
        RECT  3.070 1.345 3.300 3.700 ;
        RECT  3.300 3.625 4.225 3.965 ;
        RECT  3.030 0.630 5.630 0.970 ;
        RECT  1.825 0.885 3.370 1.115 ;
        RECT  1.825 0.885 2.110 1.450 ;
        RECT  5.990 0.980 6.330 1.850 ;
        RECT  5.780 1.620 7.290 1.850 ;
        RECT  6.950 1.620 7.290 1.960 ;
        RECT  5.780 1.620 6.010 2.935 ;
        RECT  4.235 2.595 6.010 2.935 ;
        RECT  7.430 0.980 7.770 1.320 ;
        RECT  4.495 1.805 4.835 2.145 ;
        RECT  3.775 1.915 4.835 2.145 ;
        RECT  3.530 2.740 4.005 3.080 ;
        RECT  3.775 1.915 4.005 3.395 ;
        RECT  3.775 3.165 7.770 3.395 ;
        RECT  7.535 0.980 7.770 3.550 ;
        RECT  7.190 2.645 7.770 3.550 ;
        RECT  12.045 2.075 12.580 2.415 ;
        RECT  8.690 1.240 9.030 3.910 ;
        RECT  12.045 2.075 12.275 3.910 ;
        RECT  8.690 3.680 12.275 3.910 ;
        RECT  0.965 3.470 2.30 3.700 ;
        RECT  3.030 0.630 4.20 0.970 ;
        RECT  3.775 3.165 6.80 3.395 ;
        RECT  8.690 3.680 11.60 3.910 ;
    END
END DLHRSX4

MACRO DLHRSX2
    CLASS CORE ;
    FOREIGN DLHRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.940 1.240 9.325 3.480 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.280 2.030 2.620 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.280 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.500 1.640 5.055 2.080 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.075 1.200 2.410 ;
        RECT  0.755 1.640 1.135 2.410 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 1.240 10.600 3.480 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.190 6.805 2.635 ;
        RECT  5.765 2.190 6.805 2.420 ;
        RECT  5.765 2.080 6.105 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  8.180 -0.400 11.160 0.720 ;
        RECT  6.045 -0.400 6.385 1.320 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 4.010 11.160 5.280 ;
        RECT  8.380 4.170 9.840 5.280 ;
        RECT  6.285 3.625 6.625 5.280 ;
        RECT  4.970 3.625 5.310 5.280 ;
        RECT  1.540 3.930 2.900 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.795 ;
        RECT  1.365 1.565 2.245 1.795 ;
        RECT  1.960 1.565 2.245 1.905 ;
        RECT  0.180 0.630 0.410 2.870 ;
        RECT  0.180 2.640 1.080 2.870 ;
        RECT  0.740 2.640 1.080 3.150 ;
        RECT  2.475 1.090 3.340 1.335 ;
        RECT  0.170 3.100 0.510 3.610 ;
        RECT  2.475 1.090 2.705 3.700 ;
        RECT  1.995 2.850 2.705 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 4.080 3.700 ;
        RECT  3.740 3.470 4.080 4.010 ;
        RECT  1.775 0.630 4.770 0.860 ;
        RECT  1.775 0.630 2.110 1.035 ;
        RECT  1.785 0.630 2.110 1.045 ;
        RECT  4.430 0.630 4.770 1.310 ;
        RECT  5.285 0.980 5.665 1.850 ;
        RECT  2.935 1.565 3.220 1.905 ;
        RECT  5.285 1.620 6.905 1.850 ;
        RECT  2.935 1.675 4.250 1.905 ;
        RECT  6.565 1.620 6.905 1.960 ;
        RECT  4.020 1.675 4.250 2.630 ;
        RECT  4.020 2.290 4.360 2.630 ;
        RECT  4.020 2.400 5.515 2.630 ;
        RECT  5.285 0.980 5.515 2.935 ;
        RECT  5.285 2.650 5.865 2.935 ;
        RECT  6.805 0.980 7.385 1.320 ;
        RECT  3.350 2.180 3.690 2.520 ;
        RECT  3.460 2.180 3.690 3.240 ;
        RECT  7.045 2.645 7.385 3.395 ;
        RECT  3.460 3.010 4.890 3.240 ;
        RECT  7.150 0.980 7.385 3.395 ;
        RECT  4.660 3.165 7.385 3.395 ;
        RECT  7.620 1.170 7.960 3.940 ;
        RECT  7.620 3.710 10.410 3.940 ;
        RECT  10.070 3.710 10.410 4.070 ;
        RECT  0.965 3.470 3.40 3.700 ;
        RECT  1.775 0.630 3.90 0.860 ;
        RECT  4.660 3.165 6.40 3.395 ;
        RECT  7.620 3.710 9.60 3.940 ;
    END
END DLHRSX2

MACRO DLHRSX1
    CLASS CORE ;
    FOREIGN DLHRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.860 2.250 9.325 2.630 ;
        RECT  8.750 3.270 9.090 4.180 ;
        RECT  8.860 1.220 9.090 4.180 ;
        RECT  8.750 1.220 9.090 1.560 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.810 2.230 2.400 2.665 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 3.270 10.585 4.180 ;
        RECT  10.190 1.240 10.530 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.285 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.400 2.070 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.075 6.805 2.635 ;
        RECT  5.995 2.075 6.805 2.320 ;
        RECT  5.995 1.975 6.335 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.585 ;
        RECT  7.950 -0.400 8.290 0.710 ;
        RECT  6.295 -0.400 6.635 1.150 ;
        RECT  1.210 -0.400 1.550 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 3.330 9.810 5.280 ;
        RECT  7.815 4.170 8.155 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.630 0.520 1.410 ;
        RECT  0.170 1.215 1.860 1.410 ;
        RECT  0.170 1.180 1.835 1.410 ;
        RECT  1.630 1.335 2.445 1.680 ;
        RECT  0.170 0.630 0.400 3.250 ;
        RECT  0.170 3.020 1.120 3.250 ;
        RECT  0.780 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 0.970 2.785 ;
        RECT  0.630 2.520 1.580 2.785 ;
        RECT  1.350 2.520 1.580 3.340 ;
        RECT  1.350 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  2.025 0.630 4.870 0.860 ;
        RECT  4.640 0.630 4.870 1.280 ;
        RECT  2.025 0.630 2.310 1.040 ;
        RECT  4.640 0.940 4.980 1.280 ;
        RECT  5.535 0.810 5.915 1.745 ;
        RECT  3.135 1.555 3.420 1.895 ;
        RECT  5.535 1.500 7.005 1.745 ;
        RECT  6.665 1.500 7.005 1.840 ;
        RECT  3.135 1.665 4.305 1.895 ;
        RECT  4.075 1.665 4.305 2.655 ;
        RECT  4.075 2.290 4.550 2.655 ;
        RECT  5.535 0.810 5.765 2.835 ;
        RECT  4.075 2.425 5.765 2.655 ;
        RECT  5.535 2.550 6.040 2.835 ;
        RECT  7.010 0.865 7.500 1.205 ;
        RECT  7.265 0.865 7.500 3.295 ;
        RECT  3.520 2.500 3.845 3.115 ;
        RECT  3.520 2.885 5.120 3.115 ;
        RECT  7.265 2.720 7.615 3.295 ;
        RECT  4.890 3.065 7.615 3.295 ;
        RECT  8.040 1.170 8.380 2.505 ;
        RECT  8.040 2.130 8.615 2.505 ;
        RECT  8.040 1.170 8.270 3.785 ;
        RECT  7.815 3.445 8.270 3.785 ;
        RECT  2.025 0.630 3.50 0.860 ;
        RECT  4.890 3.065 6.30 3.295 ;
    END
END DLHRSX1

MACRO DLHRSX0
    CLASS CORE ;
    FOREIGN DLHRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.225 2.250 8.065 2.630 ;
        RECT  7.225 0.675 7.870 1.015 ;
        RECT  6.810 3.965 7.455 4.250 ;
        RECT  7.225 0.675 7.455 4.250 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.395 2.630 ;
        RECT  1.790 2.120 2.395 2.460 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.578  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 3.795 9.335 4.135 ;
        RECT  9.105 0.630 9.335 4.135 ;
        RECT  8.930 0.630 9.335 1.410 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.090 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.270 2.280 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.560 2.230 5.900 2.755 ;
        RECT  5.165 2.230 5.900 2.630 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.225 -0.400 8.570 0.970 ;
        RECT  6.080 -0.400 6.995 1.145 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.685 3.885 8.495 5.280 ;
        RECT  5.190 3.965 6.260 5.280 ;
        RECT  1.645 3.660 2.790 5.280 ;
        RECT  0.180 3.700 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 2.395 1.410 ;
        RECT  2.055 1.180 2.395 1.790 ;
        RECT  0.115 1.200 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  0.900 3.185 1.155 4.000 ;
        RECT  0.900 3.660 1.240 4.000 ;
        RECT  2.625 1.230 3.520 1.540 ;
        RECT  0.575 2.610 0.915 2.955 ;
        RECT  0.575 2.695 1.615 2.955 ;
        RECT  2.625 1.230 2.855 3.240 ;
        RECT  1.385 2.860 2.855 3.240 ;
        RECT  1.385 3.010 3.440 3.240 ;
        RECT  3.210 3.010 3.440 4.250 ;
        RECT  3.210 3.965 4.185 4.250 ;
        RECT  1.950 0.630 2.290 0.950 ;
        RECT  1.950 0.720 4.920 0.950 ;
        RECT  4.580 0.720 4.920 1.540 ;
        RECT  5.280 1.385 5.620 2.000 ;
        RECT  3.085 1.770 6.535 2.000 ;
        RECT  3.085 1.770 3.370 2.110 ;
        RECT  6.230 1.770 6.535 2.365 ;
        RECT  4.130 1.770 4.470 2.635 ;
        RECT  6.230 1.770 6.460 3.275 ;
        RECT  5.320 2.985 6.460 3.275 ;
        RECT  3.455 2.440 3.900 2.780 ;
        RECT  3.670 2.440 3.900 3.735 ;
        RECT  6.710 3.095 6.995 3.735 ;
        RECT  6.765 1.505 6.995 3.735 ;
        RECT  3.670 3.505 6.995 3.735 ;
        RECT  7.685 1.375 8.525 1.715 ;
        RECT  8.295 2.395 8.750 2.735 ;
        RECT  8.295 1.375 8.525 3.420 ;
        RECT  7.745 3.080 8.525 3.420 ;
        RECT  0.180 1.180 1.40 1.410 ;
        RECT  1.385 3.010 2.60 3.240 ;
        RECT  1.950 0.720 3.50 0.950 ;
        RECT  3.085 1.770 5.20 2.000 ;
        RECT  3.670 3.505 5.60 3.735 ;
    END
END DLHRSX0

MACRO DLHRSQX4
    CLASS CORE ;
    FOREIGN DLHRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.140 2.030 2.480 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.140 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.065 1.640 5.545 2.145 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.214  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.200 2.420 ;
        RECT  0.755 1.640 1.135 2.420 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.450 1.130 11.845 3.880 ;
        RECT  10.170 2.130 11.845 2.360 ;
        RECT  10.010 2.640 10.400 3.880 ;
        RECT  10.170 1.130 10.400 3.880 ;
        RECT  10.010 1.130 10.400 1.470 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.240 2.250 6.805 2.635 ;
        RECT  6.240 2.080 6.570 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.730 -0.400 11.070 1.470 ;
        RECT  8.130 -0.400 9.590 0.720 ;
        RECT  6.710 -0.400 7.050 1.320 ;
        RECT  2.330 -0.400 2.670 0.655 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.730 2.640 11.070 5.280 ;
        RECT  9.250 3.950 9.590 5.280 ;
        RECT  8.000 2.640 8.310 5.280 ;
        RECT  6.430 3.625 6.770 5.280 ;
        RECT  5.185 3.900 5.525 5.280 ;
        RECT  1.540 3.930 2.920 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.910 ;
        RECT  1.365 1.680 2.730 1.910 ;
        RECT  2.500 1.680 2.730 2.610 ;
        RECT  2.510 2.290 2.840 2.625 ;
        RECT  0.180 0.630 0.410 2.880 ;
        RECT  0.180 2.650 1.080 2.880 ;
        RECT  0.740 2.650 1.080 3.150 ;
        RECT  4.060 1.235 4.400 1.575 ;
        RECT  3.070 1.345 4.400 1.575 ;
        RECT  1.995 2.740 2.310 3.700 ;
        RECT  0.170 3.110 0.510 3.610 ;
        RECT  1.995 2.775 2.335 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 3.525 3.700 ;
        RECT  0.965 3.470 2.40 3.700 ;
        RECT  3.070 1.345 3.300 3.700 ;
        RECT  3.300 3.625 4.225 3.855 ;
        RECT  3.885 3.625 4.225 3.965 ;
        RECT  3.030 0.670 5.630 0.970 ;
        RECT  5.290 0.630 5.630 0.970 ;
        RECT  1.825 0.885 3.370 1.115 ;
        RECT  1.825 0.885 2.110 1.450 ;
        RECT  5.990 0.980 6.330 1.850 ;
        RECT  5.780 1.620 7.290 1.850 ;
        RECT  6.950 1.620 7.290 1.960 ;
        RECT  5.780 1.620 6.010 2.935 ;
        RECT  4.235 2.595 6.010 2.935 ;
        RECT  7.430 0.980 7.770 1.320 ;
        RECT  4.495 1.805 4.835 2.145 ;
        RECT  3.775 1.915 4.835 2.145 ;
        RECT  3.530 2.740 4.005 3.080 ;
        RECT  3.775 1.915 4.005 3.395 ;
        RECT  3.775 3.165 7.770 3.395 ;
        RECT  7.535 0.980 7.770 3.550 ;
        RECT  7.190 2.645 7.770 3.550 ;
        RECT  8.690 2.075 9.940 2.415 ;
        RECT  8.690 1.240 9.030 3.550 ;
    END
END DLHRSQX4

MACRO DLHRSQX2
    CLASS CORE ;
    FOREIGN DLHRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 2.280 2.030 2.620 ;
        RECT  1.385 2.860 1.765 3.240 ;
        RECT  1.535 2.280 1.765 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.500 1.640 5.055 2.080 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.075 1.200 2.410 ;
        RECT  0.755 1.640 1.135 2.410 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.945 2.640 9.390 3.550 ;
        RECT  9.160 1.240 9.390 3.550 ;
        RECT  9.000 1.240 9.390 1.580 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.190 6.805 2.635 ;
        RECT  5.765 2.190 6.805 2.420 ;
        RECT  5.765 2.080 6.105 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  9.560 -0.400 9.900 0.720 ;
        RECT  8.240 -0.400 8.580 0.720 ;
        RECT  6.045 -0.400 6.385 1.320 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.560 3.950 9.900 5.280 ;
        RECT  8.440 3.950 8.780 5.280 ;
        RECT  6.285 3.625 6.625 5.280 ;
        RECT  4.970 3.625 5.310 5.280 ;
        RECT  1.540 3.930 2.900 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 1.595 1.410 ;
        RECT  1.365 1.180 1.595 1.795 ;
        RECT  1.365 1.565 2.245 1.795 ;
        RECT  1.960 1.565 2.245 1.905 ;
        RECT  0.180 0.630 0.410 2.870 ;
        RECT  0.180 2.640 1.080 2.870 ;
        RECT  0.740 2.640 1.080 3.150 ;
        RECT  2.475 1.090 3.340 1.335 ;
        RECT  0.170 3.100 0.510 3.610 ;
        RECT  2.475 1.090 2.705 3.700 ;
        RECT  1.995 2.850 2.705 3.700 ;
        RECT  0.170 3.380 1.195 3.610 ;
        RECT  0.965 3.470 4.080 3.700 ;
        RECT  3.740 3.470 4.080 4.010 ;
        RECT  1.775 0.630 4.660 0.860 ;
        RECT  4.430 0.630 4.660 1.310 ;
        RECT  1.775 0.630 2.110 1.035 ;
        RECT  1.785 0.630 2.110 1.045 ;
        RECT  4.430 0.970 4.770 1.310 ;
        RECT  5.285 0.980 5.625 1.850 ;
        RECT  2.935 1.565 3.220 1.905 ;
        RECT  5.285 1.620 6.905 1.850 ;
        RECT  2.935 1.675 4.250 1.905 ;
        RECT  6.565 1.620 6.905 1.960 ;
        RECT  4.020 1.675 4.250 2.630 ;
        RECT  4.020 2.290 4.360 2.630 ;
        RECT  4.020 2.400 5.515 2.630 ;
        RECT  5.285 0.980 5.515 2.935 ;
        RECT  5.285 2.650 5.865 2.935 ;
        RECT  6.805 0.980 7.385 1.320 ;
        RECT  3.350 2.180 3.690 2.520 ;
        RECT  3.460 2.180 3.690 3.240 ;
        RECT  7.045 2.640 7.385 3.395 ;
        RECT  3.460 3.010 4.890 3.240 ;
        RECT  7.150 0.980 7.385 3.395 ;
        RECT  4.660 3.165 7.385 3.395 ;
        RECT  7.680 1.240 8.020 1.580 ;
        RECT  7.790 2.040 8.930 2.270 ;
        RECT  8.590 2.040 8.930 2.380 ;
        RECT  7.790 1.240 8.020 3.550 ;
        RECT  7.680 3.210 8.020 3.550 ;
        RECT  0.965 3.470 3.80 3.700 ;
        RECT  1.775 0.630 3.80 0.860 ;
        RECT  4.660 3.165 6.70 3.395 ;
    END
END DLHRSQX2

MACRO DLHRSQX1
    CLASS CORE ;
    FOREIGN DLHRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.810 2.230 2.400 2.665 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.560 2.825 9.955 3.735 ;
        RECT  9.560 1.110 9.900 3.735 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.150 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.137  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.400 2.070 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.075 6.805 2.635 ;
        RECT  5.995 2.075 6.805 2.320 ;
        RECT  5.995 1.970 6.335 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.840 -0.400 9.180 1.430 ;
        RECT  6.295 -0.400 6.635 1.155 ;
        RECT  1.210 -0.400 1.550 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.840 2.885 9.180 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.630 0.520 1.410 ;
        RECT  0.170 1.210 1.860 1.410 ;
        RECT  0.170 1.180 1.835 1.410 ;
        RECT  1.630 1.335 2.445 1.680 ;
        RECT  0.170 0.630 0.400 3.250 ;
        RECT  0.170 3.020 1.120 3.250 ;
        RECT  0.780 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 0.970 2.785 ;
        RECT  0.630 2.520 1.580 2.785 ;
        RECT  1.350 2.520 1.580 3.340 ;
        RECT  1.350 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  2.000 0.630 4.870 0.860 ;
        RECT  4.640 0.630 4.870 1.280 ;
        RECT  2.000 0.630 2.310 1.015 ;
        RECT  2.025 0.630 2.310 1.040 ;
        RECT  4.640 0.940 4.980 1.280 ;
        RECT  5.535 0.845 5.915 1.740 ;
        RECT  5.535 1.500 7.005 1.740 ;
        RECT  6.665 1.500 7.005 1.840 ;
        RECT  3.135 1.555 4.305 1.895 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 4.550 2.655 ;
        RECT  4.075 2.425 5.765 2.655 ;
        RECT  5.535 0.845 5.765 2.655 ;
        RECT  5.555 2.550 6.040 2.835 ;
        RECT  7.010 0.885 7.615 1.225 ;
        RECT  3.520 2.500 3.845 3.115 ;
        RECT  3.520 2.885 5.120 3.115 ;
        RECT  7.265 0.885 7.615 3.295 ;
        RECT  4.890 3.065 7.615 3.295 ;
        RECT  7.270 0.885 7.615 3.450 ;
        RECT  8.040 0.990 8.425 1.330 ;
        RECT  8.075 1.850 9.330 2.190 ;
        RECT  8.075 0.990 8.425 3.165 ;
        RECT  2.000 0.630 3.00 0.860 ;
        RECT  4.890 3.065 6.60 3.295 ;
    END
END DLHRSQX1

MACRO DLHRSQX0
    CLASS CORE ;
    FOREIGN DLHRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.120 2.395 2.630 ;
        RECT  1.790 2.120 2.395 2.460 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.185 2.995 8.705 3.335 ;
        RECT  8.475 1.360 8.705 3.335 ;
        RECT  8.295 1.360 8.705 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.090 3.275 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.270 2.280 ;
        END
    END SN
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.560 2.230 5.900 2.755 ;
        RECT  5.165 2.230 5.900 2.630 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  8.225 -0.400 8.570 0.900 ;
        RECT  6.080 -0.400 6.995 1.145 ;
        RECT  1.010 -0.400 1.350 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.685 3.795 8.470 5.280 ;
        RECT  5.080 3.965 6.260 5.280 ;
        RECT  1.645 3.660 2.790 5.280 ;
        RECT  0.180 3.700 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 1.410 ;
        RECT  0.180 1.180 2.395 1.410 ;
        RECT  2.055 1.180 2.395 1.790 ;
        RECT  0.115 1.200 0.345 3.470 ;
        RECT  0.115 3.185 1.155 3.470 ;
        RECT  0.900 3.185 1.155 4.000 ;
        RECT  0.900 3.660 1.240 4.000 ;
        RECT  2.625 1.230 3.520 1.540 ;
        RECT  0.575 2.610 0.915 2.955 ;
        RECT  0.575 2.695 1.615 2.955 ;
        RECT  2.625 1.230 2.855 3.240 ;
        RECT  1.385 2.860 2.855 3.240 ;
        RECT  1.385 3.010 3.440 3.240 ;
        RECT  3.210 3.010 3.440 4.250 ;
        RECT  3.210 3.965 4.185 4.250 ;
        RECT  1.950 0.630 2.290 0.950 ;
        RECT  1.950 0.720 4.920 0.950 ;
        RECT  4.580 0.720 4.920 1.540 ;
        RECT  5.280 1.385 5.620 2.000 ;
        RECT  3.085 1.770 6.535 2.000 ;
        RECT  3.085 1.770 3.370 2.110 ;
        RECT  6.230 1.770 6.535 2.365 ;
        RECT  4.130 1.770 4.470 2.635 ;
        RECT  6.230 1.770 6.460 3.275 ;
        RECT  5.320 2.985 6.460 3.275 ;
        RECT  3.455 2.440 3.900 2.780 ;
        RECT  3.670 2.440 3.900 3.735 ;
        RECT  6.710 3.095 6.995 3.735 ;
        RECT  6.765 1.505 6.995 3.735 ;
        RECT  3.670 3.505 6.995 3.735 ;
        RECT  7.510 0.655 7.850 2.615 ;
        RECT  7.225 2.275 8.155 2.615 ;
        RECT  7.225 2.275 7.455 4.250 ;
        RECT  6.860 3.965 7.455 4.250 ;
        RECT  0.180 1.180 1.50 1.410 ;
        RECT  1.385 3.010 2.60 3.240 ;
        RECT  1.950 0.720 3.60 0.950 ;
        RECT  3.085 1.770 5.30 2.000 ;
        RECT  3.670 3.505 5.20 3.735 ;
    END
END DLHRSQX0

MACRO DLHRQX4
    CLASS CORE ;
    FOREIGN DLHRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.383  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.900 3.025 6.280 3.385 ;
        RECT  5.780 2.855 6.235 3.260 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.190 1.130 10.585 3.880 ;
        RECT  8.750 2.180 10.585 2.410 ;
        RECT  8.750 1.130 9.090 3.880 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.190 1.670 2.420 ;
        RECT  1.330 2.080 1.670 2.420 ;
        RECT  0.755 2.190 1.135 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.470 ;
        RECT  6.870 -0.400 8.330 0.720 ;
        RECT  5.450 -0.400 5.790 1.205 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.470 2.640 9.810 5.280 ;
        RECT  7.990 3.950 8.330 5.280 ;
        RECT  6.670 2.925 7.010 5.280 ;
        RECT  4.545 4.150 4.885 5.280 ;
        RECT  2.205 3.900 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  3.875 2.455 4.215 2.795 ;
        RECT  0.180 2.645 0.520 3.460 ;
        RECT  3.875 2.455 4.105 3.460 ;
        RECT  0.180 3.230 4.105 3.460 ;
        RECT  1.700 0.980 2.130 1.850 ;
        RECT  0.660 1.620 2.130 1.850 ;
        RECT  0.660 1.620 1.000 1.960 ;
        RECT  3.940 1.785 4.225 2.125 ;
        RECT  3.315 1.895 4.225 2.125 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.660 2.130 3.000 ;
        RECT  3.315 1.895 3.545 3.000 ;
        RECT  1.700 2.700 3.545 3.000 ;
        RECT  2.460 0.630 2.800 0.955 ;
        RECT  4.690 0.630 5.145 0.955 ;
        RECT  2.460 0.725 5.145 0.955 ;
        RECT  4.915 0.630 5.145 1.665 ;
        RECT  6.170 1.085 6.510 1.665 ;
        RECT  4.915 1.435 6.510 1.665 ;
        RECT  3.660 1.215 4.000 1.555 ;
        RECT  3.660 1.325 4.685 1.555 ;
        RECT  4.455 1.895 7.200 2.125 ;
        RECT  6.860 1.895 7.200 2.235 ;
        RECT  4.455 1.325 4.685 3.920 ;
        RECT  5.345 3.470 5.685 3.920 ;
        RECT  3.435 3.690 5.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  4.915 2.355 6.630 2.585 ;
        RECT  4.915 2.355 5.200 2.695 ;
        RECT  6.410 2.465 7.770 2.695 ;
        RECT  7.430 1.240 7.770 3.550 ;
        RECT  0.180 3.230 3.40 3.460 ;
        RECT  2.460 0.725 4.80 0.955 ;
        RECT  4.455 1.895 6.40 2.125 ;
        RECT  3.435 3.690 4.90 3.920 ;
    END
END DLHRQX4

MACRO DLHRQX2
    CLASS CORE ;
    FOREIGN DLHRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.140 2.595 3.655 3.240 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.755 1.640 6.315 2.085 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.240 1.140 3.550 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 2.190 8.065 2.635 ;
        RECT  7.150 2.190 8.065 2.420 ;
        RECT  7.150 2.080 7.490 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.540 -0.400 7.880 1.320 ;
        RECT  2.620 -0.400 2.960 0.765 ;
        RECT  1.560 -0.400 1.900 0.720 ;
        RECT  0.240 -0.400 0.580 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.540 3.680 7.880 5.280 ;
        RECT  6.225 3.680 6.565 5.280 ;
        RECT  3.935 3.930 4.275 5.280 ;
        RECT  1.360 3.950 1.700 5.280 ;
        RECT  0.240 3.950 0.580 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.010 1.240 2.460 1.795 ;
        RECT  2.010 1.565 3.855 1.795 ;
        RECT  3.570 1.565 3.855 1.905 ;
        RECT  2.010 1.240 2.240 3.550 ;
        RECT  2.010 2.640 2.460 3.550 ;
        RECT  4.085 1.090 4.950 1.335 ;
        RECT  2.470 2.025 2.810 2.365 ;
        RECT  2.470 2.135 4.315 2.365 ;
        RECT  4.085 1.090 4.315 3.700 ;
        RECT  3.135 3.470 5.335 3.700 ;
        RECT  3.135 3.470 3.475 3.810 ;
        RECT  4.995 3.470 5.335 3.810 ;
        RECT  3.380 0.630 6.380 0.860 ;
        RECT  3.380 0.630 3.720 1.215 ;
        RECT  6.040 0.630 6.380 1.310 ;
        RECT  6.690 0.980 7.120 1.850 ;
        RECT  4.545 1.565 4.830 1.905 ;
        RECT  6.690 1.620 8.160 1.850 ;
        RECT  4.545 1.675 5.505 1.905 ;
        RECT  7.820 1.620 8.160 1.960 ;
        RECT  5.275 1.675 5.505 2.780 ;
        RECT  6.690 0.980 6.920 2.990 ;
        RECT  5.275 2.480 6.920 2.780 ;
        RECT  6.690 2.650 7.120 2.990 ;
        RECT  8.300 0.980 8.640 1.320 ;
        RECT  4.605 2.235 4.945 2.575 ;
        RECT  4.715 2.235 4.945 3.240 ;
        RECT  4.715 3.010 6.145 3.240 ;
        RECT  5.915 3.220 8.640 3.450 ;
        RECT  8.405 0.980 8.640 3.455 ;
        RECT  8.300 2.645 8.640 3.455 ;
        RECT  3.135 3.470 4.50 3.700 ;
        RECT  3.380 0.630 5.60 0.860 ;
        RECT  5.915 3.220 7.80 3.450 ;
    END
END DLHRQX2

MACRO DLHRQX1
    CLASS CORE ;
    FOREIGN DLHRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.176  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.480 1.615 3.035 2.060 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 2.970 1.240 3.880 ;
        RECT  0.900 0.700 1.240 1.040 ;
        RECT  0.900 0.700 1.135 3.880 ;
        RECT  0.755 2.250 1.135 2.630 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.840 2.095 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 2.075 7.435 2.635 ;
        RECT  6.570 2.075 7.435 2.320 ;
        RECT  6.570 1.980 6.855 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.945 -0.400 7.285 1.270 ;
        RECT  2.135 -0.400 2.475 0.710 ;
        RECT  0.180 -0.400 0.520 1.060 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.910 3.525 7.250 5.280 ;
        RECT  5.810 3.800 6.150 5.280 ;
        RECT  2.465 3.530 3.500 5.280 ;
        RECT  0.180 2.960 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.530 1.360 1.870 1.700 ;
        RECT  1.530 1.360 1.795 2.755 ;
        RECT  1.365 2.415 1.795 2.755 ;
        RECT  1.565 1.360 1.795 3.850 ;
        RECT  1.565 3.510 2.085 3.850 ;
        RECT  4.125 1.090 4.465 1.375 ;
        RECT  3.440 1.145 4.465 1.375 ;
        RECT  2.025 2.440 2.325 3.050 ;
        RECT  3.440 1.145 3.670 3.050 ;
        RECT  2.025 2.710 3.670 3.050 ;
        RECT  2.025 2.750 3.960 3.050 ;
        RECT  3.730 2.750 3.960 3.830 ;
        RECT  3.730 3.600 4.790 3.830 ;
        RECT  4.450 3.600 4.790 3.940 ;
        RECT  2.895 0.630 5.865 0.860 ;
        RECT  2.895 0.630 3.235 1.040 ;
        RECT  5.525 0.630 5.865 1.375 ;
        RECT  6.225 0.810 6.565 1.730 ;
        RECT  6.110 1.500 7.530 1.730 ;
        RECT  7.190 1.500 7.530 1.840 ;
        RECT  3.900 1.605 4.915 1.945 ;
        RECT  4.685 1.605 4.915 2.835 ;
        RECT  6.110 1.495 6.340 2.835 ;
        RECT  4.685 2.415 6.340 2.835 ;
        RECT  4.685 2.550 6.435 2.835 ;
        RECT  7.665 0.865 8.010 1.205 ;
        RECT  7.660 2.820 8.010 3.295 ;
        RECT  7.775 0.865 8.010 3.295 ;
        RECT  4.190 3.065 8.010 3.295 ;
        RECT  4.190 3.010 4.530 3.350 ;
        RECT  2.895 0.630 4.50 0.860 ;
        RECT  4.190 3.065 7.70 3.295 ;
    END
END DLHRQX1

MACRO DLHRQX0
    CLASS CORE ;
    FOREIGN DLHRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.230 6.245 2.755 ;
        END
    END G
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.640 2.110 2.110 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.350 0.660 1.160 1.000 ;
        RECT  0.125 2.800 0.795 3.240 ;
        RECT  0.350 0.660 0.580 3.240 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.860 5.345 3.240 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.310 -0.400 6.650 1.120 ;
        RECT  1.680 -0.400 2.020 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  5.410 3.965 6.590 5.280 ;
        RECT  1.955 3.660 3.120 5.280 ;
        RECT  0.455 3.600 0.795 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.810 1.360 1.150 2.570 ;
        RECT  2.440 2.200 2.725 2.570 ;
        RECT  0.810 2.340 2.725 2.570 ;
        RECT  1.025 2.340 1.255 4.000 ;
        RECT  1.025 3.660 1.495 4.000 ;
        RECT  2.955 1.200 3.850 1.540 ;
        RECT  2.955 1.200 3.185 3.240 ;
        RECT  2.385 2.860 3.185 3.240 ;
        RECT  1.485 3.010 3.770 3.240 ;
        RECT  1.485 3.010 1.775 3.420 ;
        RECT  3.540 3.010 3.770 4.250 ;
        RECT  3.540 3.965 4.395 4.250 ;
        RECT  2.480 0.630 2.820 0.970 ;
        RECT  2.480 0.740 5.250 0.970 ;
        RECT  4.910 0.740 5.250 1.540 ;
        RECT  5.610 1.360 5.950 2.000 ;
        RECT  3.415 1.770 6.865 2.000 ;
        RECT  3.415 1.770 4.800 2.110 ;
        RECT  6.560 1.770 6.865 2.365 ;
        RECT  4.460 1.770 4.800 2.540 ;
        RECT  6.560 1.770 6.790 3.275 ;
        RECT  5.650 2.985 6.790 3.275 ;
        RECT  7.070 1.360 7.380 1.665 ;
        RECT  3.785 2.440 4.230 2.780 ;
        RECT  4.000 2.440 4.230 3.735 ;
        RECT  7.040 3.140 7.380 3.735 ;
        RECT  7.095 1.360 7.380 3.735 ;
        RECT  4.000 3.505 7.380 3.735 ;
        RECT  1.485 3.010 2.70 3.240 ;
        RECT  2.480 0.740 4.30 0.970 ;
        RECT  3.415 1.770 5.20 2.000 ;
        RECT  4.000 3.505 6.60 3.735 ;
    END
END DLHRQX0

MACRO DLHQX4
    CLASS CORE ;
    FOREIGN DLHQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.485 1.640 3.035 2.125 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 1.130 8.695 3.880 ;
        RECT  6.860 2.180 8.695 2.410 ;
        RECT  6.860 1.130 7.200 3.880 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.190 1.670 2.420 ;
        RECT  1.330 2.080 1.670 2.420 ;
        RECT  0.755 2.190 1.135 2.635 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.470 ;
        RECT  6.100 -0.400 6.440 0.720 ;
        RECT  4.780 -0.400 5.120 0.985 ;
        RECT  2.460 -0.400 2.800 0.955 ;
        RECT  0.940 -0.400 1.280 1.320 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 2.640 7.920 5.280 ;
        RECT  6.100 2.910 6.440 5.280 ;
        RECT  4.545 4.150 4.885 5.280 ;
        RECT  2.205 3.785 2.545 5.280 ;
        RECT  0.940 3.690 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.980 0.520 1.320 ;
        RECT  0.180 0.980 0.415 3.460 ;
        RECT  0.180 2.645 0.520 3.460 ;
        RECT  3.875 2.455 4.215 3.460 ;
        RECT  0.180 3.230 4.215 3.460 ;
        RECT  1.700 0.980 2.130 1.850 ;
        RECT  0.660 1.620 2.130 1.850 ;
        RECT  0.660 1.620 1.000 1.960 ;
        RECT  3.940 1.785 4.225 2.125 ;
        RECT  3.315 1.895 4.225 2.125 ;
        RECT  1.900 0.980 2.130 3.000 ;
        RECT  1.700 2.660 2.130 3.000 ;
        RECT  3.315 1.895 3.545 3.000 ;
        RECT  1.700 2.700 3.545 3.000 ;
        RECT  3.660 1.215 4.000 1.555 ;
        RECT  3.660 1.325 4.685 1.555 ;
        RECT  4.455 1.860 6.120 2.090 ;
        RECT  5.780 1.860 6.120 2.220 ;
        RECT  4.455 1.325 4.685 3.920 ;
        RECT  3.435 3.690 4.685 3.920 ;
        RECT  3.435 3.690 3.775 4.030 ;
        RECT  5.540 1.240 6.580 1.580 ;
        RECT  4.915 2.320 5.235 2.680 ;
        RECT  6.350 1.240 6.580 2.680 ;
        RECT  4.915 2.450 6.580 2.680 ;
        RECT  5.305 2.450 5.645 4.170 ;
        RECT  0.180 3.230 3.80 3.460 ;
    END
END DLHQX4

MACRO DLHQX2
    CLASS CORE ;
    FOREIGN DLHQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.615 5.160 2.080 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.240 1.140 3.550 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.190 6.805 2.635 ;
        RECT  5.890 2.190 6.805 2.420 ;
        RECT  5.890 2.080 6.230 2.420 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.320 ;
        RECT  4.900 -0.400 5.240 0.850 ;
        RECT  2.930 -0.400 3.270 0.810 ;
        RECT  1.560 -0.400 1.900 0.720 ;
        RECT  0.240 -0.400 0.580 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.480 3.950 6.820 5.280 ;
        RECT  5.110 3.750 5.450 5.280 ;
        RECT  2.560 3.910 2.905 5.280 ;
        RECT  1.360 3.950 1.700 5.280 ;
        RECT  0.240 3.950 0.580 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.930 1.240 2.460 1.580 ;
        RECT  1.930 1.240 2.160 3.550 ;
        RECT  1.930 2.690 2.785 3.030 ;
        RECT  1.930 2.690 2.460 3.550 ;
        RECT  3.855 0.630 4.195 1.415 ;
        RECT  3.015 1.180 4.195 1.415 ;
        RECT  2.390 2.020 3.245 2.360 ;
        RECT  3.015 1.180 3.245 3.190 ;
        RECT  3.135 2.970 3.365 4.035 ;
        RECT  3.135 3.750 4.220 4.035 ;
        RECT  5.600 0.980 5.940 1.850 ;
        RECT  5.430 1.620 6.900 1.850 ;
        RECT  6.560 1.620 6.900 1.960 ;
        RECT  3.575 1.680 4.295 2.020 ;
        RECT  5.430 1.620 5.660 3.060 ;
        RECT  4.065 1.680 4.295 3.060 ;
        RECT  4.065 2.720 4.500 3.060 ;
        RECT  5.430 2.650 5.990 3.060 ;
        RECT  4.065 2.830 5.990 3.060 ;
        RECT  7.040 0.980 7.380 1.320 ;
        RECT  3.490 2.350 3.830 2.690 ;
        RECT  3.600 2.350 3.830 3.520 ;
        RECT  7.040 2.645 7.380 3.520 ;
        RECT  7.145 0.980 7.380 3.520 ;
        RECT  3.600 3.290 7.380 3.520 ;
        RECT  3.600 3.290 6.90 3.520 ;
    END
END DLHQX2

MACRO DLHQX1
    CLASS CORE ;
    FOREIGN DLHQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.758  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.945 0.700 1.285 3.880 ;
        RECT  0.755 2.250 1.285 2.630 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.210 2.095 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.075 6.805 2.635 ;
        RECT  5.940 2.075 6.805 2.320 ;
        RECT  5.940 1.980 6.225 2.320 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.315 -0.400 6.655 1.270 ;
        RECT  4.895 -0.400 5.235 1.375 ;
        RECT  1.795 -0.400 2.605 0.710 ;
        RECT  0.220 -0.400 0.565 1.125 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.280 3.525 6.620 5.280 ;
        RECT  5.180 3.800 5.520 5.280 ;
        RECT  2.465 3.530 2.870 5.280 ;
        RECT  0.220 2.970 0.565 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.515 1.360 1.870 1.700 ;
        RECT  1.515 1.360 1.795 3.850 ;
        RECT  1.515 2.940 1.805 3.850 ;
        RECT  1.515 3.510 2.085 3.850 ;
        RECT  3.495 1.035 3.835 1.375 ;
        RECT  2.810 1.145 3.835 1.375 ;
        RECT  2.810 1.145 3.040 2.545 ;
        RECT  2.025 2.205 3.040 2.545 ;
        RECT  2.025 2.245 3.330 2.545 ;
        RECT  3.100 2.245 3.330 3.830 ;
        RECT  3.100 3.600 4.160 3.830 ;
        RECT  3.820 3.600 4.160 3.940 ;
        RECT  5.595 0.810 5.935 1.730 ;
        RECT  5.480 1.500 6.900 1.730 ;
        RECT  6.560 1.500 6.900 1.840 ;
        RECT  3.270 1.605 4.285 1.945 ;
        RECT  4.055 1.605 4.285 2.835 ;
        RECT  4.055 2.415 4.570 2.835 ;
        RECT  5.480 1.495 5.710 2.835 ;
        RECT  4.055 2.550 5.805 2.835 ;
        RECT  7.035 0.865 7.380 1.205 ;
        RECT  7.030 2.820 7.380 3.295 ;
        RECT  7.145 0.865 7.380 3.295 ;
        RECT  3.560 3.065 7.380 3.295 ;
        RECT  3.560 3.010 3.900 3.350 ;
        RECT  3.560 3.065 6.50 3.295 ;
    END
END DLHQX1

MACRO DLHQX0
    CLASS CORE ;
    FOREIGN DLHQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.015 0.815 3.380 ;
        RECT  0.125 2.860 0.720 3.380 ;
        RECT  0.380 1.360 0.720 3.380 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.860 4.715 3.240 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.150 2.230 5.615 2.755 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.680 -0.400 6.020 1.090 ;
        RECT  4.280 -0.400 4.620 1.540 ;
        RECT  1.980 -0.400 2.320 0.980 ;
        RECT  0.380 -0.400 0.720 0.900 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  4.780 3.965 5.960 5.280 ;
        RECT  2.175 3.470 2.515 5.280 ;
        RECT  0.475 3.930 0.815 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.180 1.250 1.520 2.540 ;
        RECT  1.180 2.200 2.095 2.540 ;
        RECT  1.050 2.310 1.280 4.160 ;
        RECT  1.050 3.890 1.615 4.160 ;
        RECT  2.880 0.640 3.220 1.540 ;
        RECT  2.325 1.310 3.220 1.540 ;
        RECT  2.325 1.310 2.555 3.240 ;
        RECT  1.510 3.010 3.140 3.240 ;
        RECT  1.510 3.010 1.850 3.365 ;
        RECT  2.910 3.010 3.140 4.250 ;
        RECT  2.910 3.965 3.650 4.250 ;
        RECT  4.980 1.360 5.320 2.000 ;
        RECT  2.785 1.770 6.235 2.000 ;
        RECT  2.785 1.770 4.170 2.110 ;
        RECT  5.930 1.770 6.235 2.365 ;
        RECT  3.830 1.770 4.170 2.540 ;
        RECT  5.930 1.770 6.160 3.275 ;
        RECT  5.020 2.985 6.160 3.275 ;
        RECT  6.440 1.360 6.750 1.665 ;
        RECT  3.155 2.440 3.600 2.780 ;
        RECT  3.370 2.440 3.600 3.735 ;
        RECT  6.410 3.095 6.750 3.735 ;
        RECT  6.465 1.360 6.750 3.735 ;
        RECT  3.370 3.505 6.750 3.735 ;
        RECT  2.785 1.770 5.60 2.000 ;
        RECT  3.370 3.505 5.70 3.735 ;
    END
END DLHQX0

MACRO DFRX4
    CLASS CORE ;
    FOREIGN DFRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 1.130 16.885 3.770 ;
        RECT  15.170 2.250 16.885 2.630 ;
        RECT  15.170 1.130 15.510 3.935 ;
        RECT  15.050 1.130 15.510 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.078  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.565 2.860 14.890 3.240 ;
        RECT  14.660 1.700 14.890 3.240 ;
        RECT  12.170 1.700 14.890 1.930 ;
        RECT  13.610 1.130 13.950 1.930 ;
        RECT  12.565 2.860 12.945 4.180 ;
        RECT  12.565 2.640 12.930 4.180 ;
        RECT  12.170 1.130 12.510 1.930 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.550 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.770 -0.400 16.110 1.470 ;
        RECT  14.330 -0.400 14.670 1.470 ;
        RECT  12.890 -0.400 13.230 1.470 ;
        RECT  10.310 -0.400 11.090 1.160 ;
        RECT  7.700 -0.400 8.040 1.320 ;
        RECT  5.690 -0.400 6.030 0.950 ;
        RECT  1.580 -0.400 2.400 1.060 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.930 4.170 16.270 5.280 ;
        RECT  14.450 3.555 14.790 5.280 ;
        RECT  13.340 3.870 13.680 5.280 ;
        RECT  11.820 3.910 12.160 5.280 ;
        RECT  10.555 3.540 10.895 5.280 ;
        RECT  8.460 3.850 8.800 5.280 ;
        RECT  6.040 2.910 6.340 5.280 ;
        RECT  0.940 4.060 2.335 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 2.860 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.090 1.190 3.680 1.530 ;
        RECT  1.835 2.325 3.320 2.665 ;
        RECT  3.090 1.190 3.320 3.275 ;
        RECT  3.090 2.935 3.570 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  3.950 2.980 4.290 3.830 ;
        RECT  0.180 3.600 4.290 3.830 ;
        RECT  2.630 0.700 4.140 0.930 ;
        RECT  3.910 0.700 4.140 1.550 ;
        RECT  2.630 0.700 2.860 1.520 ;
        RECT  0.780 1.290 2.860 1.520 ;
        RECT  3.910 1.320 4.495 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.155 1.320 4.495 1.660 ;
        RECT  6.260 0.775 7.470 1.005 ;
        RECT  4.370 0.735 5.295 1.075 ;
        RECT  5.065 0.735 5.295 3.195 ;
        RECT  6.260 0.775 6.490 1.410 ;
        RECT  5.065 1.180 6.490 1.410 ;
        RECT  7.240 0.775 7.470 2.090 ;
        RECT  7.240 1.860 8.950 2.090 ;
        RECT  8.610 1.860 8.950 2.200 ;
        RECT  5.065 1.180 5.350 3.195 ;
        RECT  6.760 1.240 7.010 1.545 ;
        RECT  9.280 1.570 9.620 1.910 ;
        RECT  3.550 1.840 3.860 2.180 ;
        RECT  3.550 1.950 4.835 2.180 ;
        RECT  6.780 1.240 7.010 2.860 ;
        RECT  6.780 2.340 7.830 2.680 ;
        RECT  9.280 1.570 9.510 2.680 ;
        RECT  5.580 2.450 9.510 2.680 ;
        RECT  6.720 2.450 7.060 2.860 ;
        RECT  4.520 1.950 4.835 3.655 ;
        RECT  7.930 3.390 9.550 3.620 ;
        RECT  6.720 2.450 6.950 3.855 ;
        RECT  5.580 2.450 5.810 3.655 ;
        RECT  4.520 3.425 5.810 3.655 ;
        RECT  7.930 3.390 8.160 3.855 ;
        RECT  6.720 3.625 8.160 3.855 ;
        RECT  9.210 3.390 9.550 4.000 ;
        RECT  8.850 0.920 9.190 1.340 ;
        RECT  8.850 1.110 10.080 1.340 ;
        RECT  9.850 1.110 10.080 3.880 ;
        RECT  11.000 1.880 11.340 2.220 ;
        RECT  9.850 1.990 11.340 2.220 ;
        RECT  7.380 2.930 10.120 3.160 ;
        RECT  7.270 3.110 7.610 3.395 ;
        RECT  9.850 1.990 10.120 3.880 ;
        RECT  9.780 2.930 10.120 3.880 ;
        RECT  11.470 0.900 11.810 1.620 ;
        RECT  10.310 1.390 11.810 1.620 ;
        RECT  10.310 1.390 10.650 1.730 ;
        RECT  11.580 2.180 14.430 2.410 ;
        RECT  14.090 2.180 14.430 2.630 ;
        RECT  11.580 0.900 11.810 3.510 ;
        RECT  11.260 2.640 11.810 3.510 ;
        RECT  0.180 3.600 3.60 3.830 ;
        RECT  0.780 1.290 1.90 1.520 ;
        RECT  5.580 2.450 8.70 2.680 ;
        RECT  7.380 2.930 9.60 3.160 ;
        RECT  11.580 2.180 13.70 2.410 ;
    END
END DFRX4

MACRO DFRX2
    CLASS CORE ;
    FOREIGN DFRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.240 11.860 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.200 3.185 11.235 3.415 ;
        RECT  11.005 1.790 11.235 3.415 ;
        RECT  10.200 1.790 11.235 2.020 ;
        RECT  10.200 1.240 10.585 2.020 ;
        RECT  10.200 3.185 10.540 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.100 2.100 5.545 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.635 3.770 2.115 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  10.960 3.950 12.420 5.280 ;
        RECT  8.295 4.140 9.780 5.280 ;
        RECT  5.910 3.830 6.250 5.280 ;
        RECT  4.770 3.910 5.110 5.280 ;
        RECT  3.510 3.880 3.850 5.280 ;
        RECT  1.680 3.960 2.020 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.960 -0.400 12.420 0.720 ;
        RECT  9.640 -0.400 9.980 0.720 ;
        RECT  8.240 -0.400 8.580 1.060 ;
        RECT  6.650 -0.400 6.990 0.950 ;
        RECT  4.640 -0.400 4.975 0.950 ;
        RECT  3.080 -0.400 3.420 0.840 ;
        RECT  0.700 -0.400 1.040 1.010 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.700 ;
        RECT  0.115 2.640 1.455 2.870 ;
        RECT  1.115 2.640 1.455 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  2.010 0.630 2.350 0.950 ;
        RECT  1.270 0.720 2.350 0.950 ;
        RECT  1.270 0.720 1.500 2.410 ;
        RECT  1.270 2.180 1.675 2.410 ;
        RECT  1.625 2.185 1.915 2.415 ;
        RECT  0.575 3.100 0.860 3.440 ;
        RECT  1.685 2.185 1.915 3.625 ;
        RECT  0.575 3.210 1.915 3.440 ;
        RECT  1.685 3.395 2.820 3.625 ;
        RECT  2.480 3.395 2.820 3.735 ;
        RECT  4.460 1.640 5.950 1.870 ;
        RECT  5.665 1.195 5.950 1.870 ;
        RECT  4.460 1.640 4.790 2.180 ;
        RECT  5.775 2.560 6.925 2.790 ;
        RECT  6.585 2.560 6.925 2.900 ;
        RECT  2.145 2.360 2.430 3.165 ;
        RECT  2.145 2.935 3.700 3.165 ;
        RECT  3.470 2.935 3.700 3.410 ;
        RECT  5.530 2.860 6.005 3.410 ;
        RECT  5.775 1.695 6.005 3.410 ;
        RECT  3.470 3.180 6.005 3.410 ;
        RECT  5.205 0.735 6.420 0.965 ;
        RECT  6.190 0.735 6.420 1.555 ;
        RECT  5.205 0.735 5.435 1.410 ;
        RECT  3.880 1.180 5.435 1.410 ;
        RECT  3.880 1.090 4.220 1.430 ;
        RECT  6.190 1.325 7.290 1.555 ;
        RECT  1.730 1.670 2.990 1.955 ;
        RECT  7.060 1.850 7.400 2.190 ;
        RECT  7.060 1.325 7.290 2.190 ;
        RECT  2.760 1.670 2.990 2.705 ;
        RECT  2.760 2.340 3.100 2.705 ;
        RECT  4.000 1.180 4.230 2.950 ;
        RECT  2.760 2.475 4.230 2.705 ;
        RECT  4.000 2.610 4.550 2.950 ;
        RECT  7.265 1.960 7.550 3.310 ;
        RECT  7.415 0.720 8.010 1.060 ;
        RECT  8.910 2.750 9.250 3.095 ;
        RECT  7.780 2.865 9.250 3.095 ;
        RECT  7.780 0.720 8.010 3.895 ;
        RECT  7.065 3.665 8.010 3.895 ;
        RECT  7.065 3.665 7.405 4.005 ;
        RECT  8.940 0.650 9.280 2.460 ;
        RECT  8.240 2.230 9.710 2.460 ;
        RECT  9.480 2.320 10.775 2.550 ;
        RECT  8.240 2.230 8.580 2.570 ;
        RECT  10.435 2.320 10.775 2.660 ;
        RECT  9.480 2.230 9.710 3.665 ;
        RECT  8.875 3.325 9.710 3.665 ;
        RECT  3.470 3.180 5.60 3.410 ;
    END
END DFRX2

MACRO DFRX1
    CLASS CORE ;
    FOREIGN DFRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.070 1.745 3.395 2.085 ;
        RECT  3.070 1.180 3.300 2.085 ;
        RECT  2.645 1.180 3.300 1.410 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.695 2.075 5.290 2.360 ;
        RECT  4.535 2.250 4.915 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.662  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 2.250 10.585 2.630 ;
        RECT  9.640 2.870 10.435 3.100 ;
        RECT  10.205 1.320 10.435 3.100 ;
        RECT  9.490 1.320 10.435 1.550 ;
        RECT  9.380 3.325 9.870 3.610 ;
        RECT  9.640 2.870 9.870 3.610 ;
        RECT  9.490 0.700 9.720 1.550 ;
        RECT  9.380 0.700 9.720 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.820 3.270 11.215 4.180 ;
        RECT  10.820 0.820 11.160 1.160 ;
        RECT  10.820 0.820 11.050 4.180 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.100 -0.400 10.440 1.090 ;
        RECT  8.575 -0.400 8.915 1.440 ;
        RECT  6.525 -0.400 7.335 0.710 ;
        RECT  4.520 -0.400 4.860 0.925 ;
        RECT  3.060 -0.400 3.400 0.800 ;
        RECT  0.960 -0.400 1.300 0.915 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.100 3.330 10.440 5.280 ;
        RECT  8.040 4.145 8.380 5.280 ;
        RECT  5.820 3.810 6.160 5.280 ;
        RECT  4.690 3.525 5.030 5.280 ;
        RECT  3.590 3.810 3.930 5.280 ;
        RECT  1.220 4.170 1.560 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.665 0.520 0.990 ;
        RECT  0.115 2.175 1.020 2.515 ;
        RECT  0.115 0.665 0.345 3.680 ;
        RECT  0.115 3.450 0.760 3.680 ;
        RECT  0.420 3.450 0.760 3.790 ;
        RECT  1.860 0.665 2.200 0.950 ;
        RECT  1.860 0.665 2.090 1.410 ;
        RECT  1.250 1.180 2.090 1.410 ;
        RECT  0.700 2.880 1.480 3.220 ;
        RECT  1.250 1.180 1.480 3.875 ;
        RECT  1.250 3.645 2.530 3.875 ;
        RECT  2.190 3.645 2.530 3.985 ;
        RECT  5.550 1.240 5.835 1.845 ;
        RECT  4.085 1.615 5.835 1.845 ;
        RECT  4.085 1.615 4.365 2.095 ;
        RECT  4.085 1.615 4.345 2.120 ;
        RECT  5.605 1.240 5.835 2.800 ;
        RECT  6.530 2.460 6.870 2.800 ;
        RECT  5.450 2.570 6.870 2.800 ;
        RECT  1.970 2.525 2.310 3.360 ;
        RECT  5.450 2.540 5.810 3.295 ;
        RECT  3.575 3.065 5.810 3.295 ;
        RECT  1.970 3.130 3.755 3.360 ;
        RECT  5.090 0.780 6.295 1.010 ;
        RECT  3.625 1.070 4.100 1.385 ;
        RECT  5.090 0.780 5.320 1.385 ;
        RECT  3.625 1.155 5.320 1.385 ;
        RECT  6.065 0.780 6.295 1.905 ;
        RECT  1.710 1.745 2.050 2.085 ;
        RECT  6.065 1.675 7.325 1.905 ;
        RECT  6.945 1.725 7.505 2.000 ;
        RECT  1.710 1.795 2.840 2.085 ;
        RECT  2.610 1.795 2.840 2.865 ;
        RECT  2.610 2.440 3.855 2.670 ;
        RECT  3.625 1.070 3.855 2.670 ;
        RECT  3.645 2.550 4.230 2.835 ;
        RECT  2.610 2.440 2.980 2.865 ;
        RECT  7.275 1.725 7.505 3.240 ;
        RECT  7.275 2.900 7.630 3.240 ;
        RECT  7.305 1.110 7.645 1.445 ;
        RECT  7.305 1.215 7.965 1.445 ;
        RECT  7.735 1.215 7.965 2.580 ;
        RECT  7.860 2.350 8.940 2.635 ;
        RECT  7.860 2.350 8.090 3.785 ;
        RECT  7.010 3.555 8.090 3.785 ;
        RECT  7.010 3.555 7.350 3.895 ;
        RECT  8.255 1.670 8.595 2.010 ;
        RECT  8.255 1.780 9.720 2.010 ;
        RECT  9.180 1.780 9.720 2.640 ;
        RECT  9.180 2.300 9.870 2.640 ;
        RECT  9.180 1.780 9.410 3.095 ;
        RECT  8.920 2.865 9.410 3.095 ;
        RECT  8.920 2.865 9.150 4.200 ;
        RECT  8.840 3.860 9.180 4.200 ;
        RECT  3.575 3.065 4.80 3.295 ;
    END
END DFRX1

MACRO DFRX0
    CLASS CORE ;
    FOREIGN DFRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.790 3.710 9.955 3.940 ;
        RECT  9.725 0.630 9.955 3.940 ;
        RECT  9.575 3.470 9.955 3.940 ;
        RECT  9.010 0.630 9.955 0.950 ;
        RECT  8.790 3.710 9.130 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 2.220 3.655 2.685 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.000 2.135 5.545 2.630 ;
        END
    END C
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.185 1.170 10.585 2.020 ;
        RECT  10.185 3.425 10.530 3.765 ;
        RECT  10.185 1.170 10.415 3.765 ;
        END
    END QN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.590 4.170 9.930 5.280 ;
        RECT  8.040 3.230 8.325 5.280 ;
        RECT  5.300 3.630 5.640 5.280 ;
        RECT  4.420 3.910 4.760 5.280 ;
        RECT  3.490 3.910 3.830 5.280 ;
        RECT  0.780 4.100 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 0.710 ;
        RECT  8.170 -0.400 8.550 0.970 ;
        RECT  6.510 -0.400 6.795 0.970 ;
        RECT  4.560 -0.400 4.845 0.970 ;
        RECT  3.260 -0.400 3.600 0.970 ;
        RECT  0.780 -0.400 1.120 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.255 0.520 2.395 ;
        RECT  0.115 1.990 1.275 2.395 ;
        RECT  0.115 1.255 0.345 3.700 ;
        RECT  0.115 3.360 0.520 3.700 ;
        RECT  1.505 1.210 2.480 1.505 ;
        RECT  1.505 1.210 1.735 2.775 ;
        RECT  0.575 2.790 1.640 3.020 ;
        RECT  0.575 2.790 0.915 3.130 ;
        RECT  1.410 2.585 1.640 4.230 ;
        RECT  1.410 3.890 2.360 4.230 ;
        RECT  5.535 1.270 5.820 1.905 ;
        RECT  4.345 2.160 4.685 2.500 ;
        RECT  5.775 1.675 6.005 3.200 ;
        RECT  4.455 2.860 6.635 3.200 ;
        RECT  1.870 3.060 2.210 3.400 ;
        RECT  1.980 3.060 2.210 3.660 ;
        RECT  4.455 2.160 4.685 3.660 ;
        RECT  1.980 3.430 4.685 3.660 ;
        RECT  5.075 0.810 6.280 1.040 ;
        RECT  3.885 1.270 4.300 1.610 ;
        RECT  6.050 0.810 6.280 1.445 ;
        RECT  5.075 0.810 5.305 1.610 ;
        RECT  3.885 1.380 5.305 1.610 ;
        RECT  1.965 1.735 4.115 1.965 ;
        RECT  1.965 1.735 2.770 2.080 ;
        RECT  6.235 1.215 6.465 2.460 ;
        RECT  6.235 2.130 6.590 2.460 ;
        RECT  6.235 2.230 7.255 2.460 ;
        RECT  2.540 1.735 2.770 3.180 ;
        RECT  3.885 1.270 4.115 3.200 ;
        RECT  7.010 2.230 7.255 3.425 ;
        RECT  2.540 2.840 2.880 3.180 ;
        RECT  3.820 2.860 4.160 3.200 ;
        RECT  7.010 3.085 7.350 3.425 ;
        RECT  7.310 0.630 7.810 0.970 ;
        RECT  7.580 2.620 8.845 2.960 ;
        RECT  7.580 0.630 7.810 3.970 ;
        RECT  6.700 3.655 7.810 3.970 ;
        RECT  9.010 1.360 9.350 2.180 ;
        RECT  8.060 1.950 9.495 2.180 ;
        RECT  9.075 1.880 9.495 2.220 ;
        RECT  8.060 1.950 8.400 2.290 ;
        RECT  9.075 1.360 9.305 3.480 ;
        RECT  8.790 3.190 9.305 3.480 ;
        RECT  4.455 2.860 5.30 3.200 ;
        RECT  1.980 3.430 3.40 3.660 ;
        RECT  1.965 1.735 3.60 1.965 ;
    END
END DFRX0

MACRO DFRSX4
    CLASS CORE ;
    FOREIGN DFRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.085  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 1.130 17.460 3.060 ;
        RECT  15.840 2.250 17.460 2.630 ;
        RECT  15.840 2.250 16.180 3.060 ;
        RECT  15.840 1.130 16.070 3.060 ;
        RECT  15.680 1.130 16.070 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.103  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.055 2.890 15.545 3.120 ;
        RECT  15.315 1.700 15.545 3.120 ;
        RECT  12.955 1.700 15.545 1.930 ;
        RECT  13.055 2.890 14.835 3.240 ;
        RECT  14.240 1.130 14.580 1.930 ;
        RECT  13.055 2.860 13.735 3.240 ;
        RECT  13.055 2.860 13.395 4.100 ;
        RECT  12.955 0.630 13.185 1.930 ;
        RECT  12.760 0.630 13.185 0.970 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.255 1.640 11.935 2.020 ;
        RECT  11.255 1.640 11.595 2.220 ;
        END
    END SN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.420 1.660 6.965 2.105 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.470 ;
        RECT  14.960 -0.400 15.300 1.470 ;
        RECT  13.520 -0.400 13.860 1.470 ;
        RECT  10.495 -0.400 11.315 0.880 ;
        RECT  8.115 -0.400 8.455 1.320 ;
        RECT  6.105 -0.400 6.445 0.970 ;
        RECT  1.580 -0.400 2.815 0.710 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.480 3.295 16.820 5.280 ;
        RECT  15.105 3.555 15.445 5.280 ;
        RECT  13.775 3.470 14.115 5.280 ;
        RECT  12.295 4.160 12.635 5.280 ;
        RECT  11.015 3.540 11.355 5.280 ;
        RECT  8.875 3.850 9.215 5.280 ;
        RECT  6.455 2.910 6.755 5.280 ;
        RECT  2.410 3.965 2.750 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 3.275 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.505 1.190 4.095 1.530 ;
        RECT  1.835 2.325 3.735 2.665 ;
        RECT  3.505 1.190 3.735 3.275 ;
        RECT  3.505 2.935 3.985 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.705 3.735 ;
        RECT  4.365 2.980 4.705 3.735 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  3.045 0.700 4.555 0.930 ;
        RECT  4.325 0.700 4.555 1.550 ;
        RECT  3.045 0.700 3.275 1.520 ;
        RECT  0.780 1.290 3.275 1.520 ;
        RECT  4.325 1.320 4.910 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.570 1.320 4.910 1.660 ;
        RECT  6.675 0.775 7.885 1.005 ;
        RECT  4.785 0.735 5.710 1.075 ;
        RECT  5.480 0.735 5.710 3.195 ;
        RECT  6.675 0.775 6.905 1.430 ;
        RECT  5.480 1.200 6.905 1.430 ;
        RECT  7.655 0.775 7.885 2.090 ;
        RECT  7.655 1.860 9.365 2.090 ;
        RECT  9.025 1.860 9.365 2.200 ;
        RECT  5.480 1.200 5.765 3.195 ;
        RECT  7.170 1.240 7.425 1.555 ;
        RECT  9.695 1.570 10.020 1.910 ;
        RECT  3.965 1.840 4.275 2.180 ;
        RECT  3.965 1.950 5.250 2.180 ;
        RECT  7.195 1.240 7.425 2.860 ;
        RECT  7.195 2.340 8.245 2.680 ;
        RECT  9.695 1.570 9.925 2.680 ;
        RECT  5.995 2.450 9.925 2.680 ;
        RECT  7.135 2.450 7.475 2.860 ;
        RECT  4.935 1.950 5.250 3.655 ;
        RECT  8.345 3.390 9.965 3.620 ;
        RECT  7.135 2.450 7.365 3.855 ;
        RECT  5.995 2.450 6.225 3.655 ;
        RECT  4.935 3.425 6.225 3.655 ;
        RECT  8.345 3.390 8.575 3.855 ;
        RECT  7.135 3.625 8.575 3.855 ;
        RECT  9.625 3.390 9.965 4.000 ;
        RECT  9.265 0.920 9.605 1.340 ;
        RECT  9.265 1.110 10.480 1.340 ;
        RECT  10.250 1.110 10.480 3.880 ;
        RECT  11.925 2.370 12.265 2.710 ;
        RECT  10.250 2.480 12.265 2.710 ;
        RECT  7.795 2.930 10.535 3.160 ;
        RECT  7.685 3.110 8.025 3.395 ;
        RECT  10.250 2.480 10.535 3.880 ;
        RECT  10.195 2.930 10.535 3.880 ;
        RECT  10.710 1.140 12.505 1.370 ;
        RECT  10.710 1.140 10.995 1.480 ;
        RECT  12.165 1.140 12.505 1.620 ;
        RECT  12.495 2.310 15.085 2.540 ;
        RECT  14.745 2.310 15.085 2.650 ;
        RECT  12.495 1.390 12.725 3.170 ;
        RECT  11.735 2.940 12.725 3.170 ;
        RECT  11.735 2.940 12.075 3.760 ;
        RECT  2.030 3.505 3.70 3.735 ;
        RECT  0.180 3.600 1.60 3.830 ;
        RECT  0.780 1.290 2.60 1.520 ;
        RECT  5.995 2.450 8.90 2.680 ;
        RECT  10.250 2.480 11.70 2.710 ;
        RECT  7.795 2.930 9.00 3.160 ;
        RECT  12.495 2.310 14.30 2.540 ;
    END
END DFRSX4

MACRO DFRSX2
    CLASS CORE ;
    FOREIGN DFRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 1.240 13.120 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.899  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.460 2.860 12.495 3.090 ;
        RECT  12.265 1.180 12.495 3.090 ;
        RECT  11.460 1.180 12.495 1.410 ;
        RECT  11.460 0.840 11.845 1.410 ;
        RECT  11.460 2.860 11.800 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.760 2.075 6.175 2.660 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.800 2.250 10.585 2.705 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 1.630 4.400 2.110 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.220 3.950 13.680 5.280 ;
        RECT  10.715 3.940 11.055 5.280 ;
        RECT  9.235 3.865 9.575 5.280 ;
        RECT  6.940 3.470 7.280 5.280 ;
        RECT  5.640 3.525 5.980 5.280 ;
        RECT  4.340 3.525 4.680 5.280 ;
        RECT  1.700 3.910 2.550 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.220 -0.400 13.680 0.720 ;
        RECT  10.740 -0.400 11.080 1.060 ;
        RECT  9.205 -0.400 9.545 1.090 ;
        RECT  7.280 -0.400 7.620 0.890 ;
        RECT  5.270 -0.400 5.610 0.925 ;
        RECT  3.640 -0.400 3.980 0.725 ;
        RECT  1.130 -0.400 1.470 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.700 ;
        RECT  0.115 2.585 2.040 2.815 ;
        RECT  1.730 2.585 2.040 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  1.700 1.035 2.780 1.325 ;
        RECT  1.700 1.035 1.930 2.355 ;
        RECT  1.700 2.125 2.500 2.355 ;
        RECT  0.575 3.100 0.915 3.440 ;
        RECT  2.270 2.125 2.500 3.575 ;
        RECT  0.575 3.210 2.500 3.440 ;
        RECT  2.270 3.345 3.350 3.575 ;
        RECT  3.010 3.345 3.350 3.685 ;
        RECT  6.300 1.240 6.590 1.845 ;
        RECT  5.090 1.615 6.635 1.845 ;
        RECT  5.090 1.615 5.430 2.100 ;
        RECT  6.405 1.615 6.635 3.295 ;
        RECT  6.405 2.280 8.035 2.510 ;
        RECT  7.695 2.280 8.035 2.605 ;
        RECT  2.730 2.310 3.060 2.650 ;
        RECT  2.830 2.310 3.060 3.115 ;
        RECT  6.400 2.780 6.740 3.295 ;
        RECT  2.830 2.885 4.330 3.115 ;
        RECT  6.405 2.280 6.740 3.295 ;
        RECT  4.100 3.065 6.740 3.295 ;
        RECT  5.840 0.780 7.050 1.010 ;
        RECT  6.820 0.780 7.050 1.390 ;
        RECT  5.840 0.780 6.070 1.385 ;
        RECT  4.510 1.155 6.070 1.385 ;
        RECT  6.820 1.160 7.435 1.390 ;
        RECT  4.510 1.070 4.850 1.410 ;
        RECT  2.160 1.555 2.500 1.895 ;
        RECT  7.205 1.160 7.435 2.010 ;
        RECT  7.205 1.670 7.545 2.010 ;
        RECT  2.160 1.665 3.620 1.895 ;
        RECT  7.205 1.780 8.495 2.010 ;
        RECT  3.390 1.665 3.620 2.655 ;
        RECT  3.390 2.290 3.730 2.655 ;
        RECT  4.630 1.155 4.860 2.835 ;
        RECT  3.390 2.425 4.860 2.655 ;
        RECT  4.630 2.550 5.220 2.835 ;
        RECT  8.265 1.780 8.495 3.065 ;
        RECT  7.635 2.835 8.495 3.065 ;
        RECT  7.635 2.835 7.865 4.040 ;
        RECT  7.635 3.810 8.795 4.040 ;
        RECT  8.485 3.805 8.795 4.100 ;
        RECT  8.455 3.810 8.795 4.100 ;
        RECT  8.175 0.630 8.955 0.950 ;
        RECT  8.725 2.965 10.720 3.250 ;
        RECT  8.725 0.630 8.955 3.525 ;
        RECT  8.095 3.295 8.955 3.525 ;
        RECT  8.095 3.295 8.435 3.580 ;
        RECT  10.540 1.560 10.880 2.020 ;
        RECT  9.185 1.790 11.180 2.020 ;
        RECT  10.950 2.120 12.035 2.460 ;
        RECT  9.185 1.790 9.470 2.700 ;
        RECT  10.950 1.790 11.180 3.710 ;
        RECT  9.965 3.480 11.180 3.710 ;
        RECT  9.965 3.480 10.305 4.070 ;
        RECT  4.100 3.065 5.20 3.295 ;
    END
END DFRSX2

MACRO DFRSX1
    CLASS CORE ;
    FOREIGN DFRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.230 1.640 4.570 2.085 ;
        RECT  3.905 1.640 4.570 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.955 2.075 6.415 2.360 ;
        RECT  5.795 2.250 6.175 2.635 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.640 10.585 2.305 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 2.250 12.475 2.630 ;
        RECT  11.530 2.870 12.325 3.100 ;
        RECT  12.095 1.235 12.325 3.100 ;
        RECT  11.380 1.235 12.325 1.465 ;
        RECT  11.270 3.665 11.760 4.005 ;
        RECT  11.530 2.870 11.760 4.005 ;
        RECT  11.380 0.700 11.610 1.465 ;
        RECT  11.270 0.700 11.610 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 0.820 13.105 4.180 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.990 -0.400 12.330 1.005 ;
        RECT  10.015 -0.400 10.355 0.880 ;
        RECT  7.725 -0.400 8.065 0.820 ;
        RECT  5.665 -0.400 6.005 0.925 ;
        RECT  4.165 -0.400 4.505 1.410 ;
        RECT  1.340 -0.400 1.680 1.565 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  11.990 3.330 12.330 5.280 ;
        RECT  10.570 4.005 10.910 5.280 ;
        RECT  9.210 3.910 9.550 5.280 ;
        RECT  7.110 3.320 7.450 5.280 ;
        RECT  5.810 3.525 6.150 5.280 ;
        RECT  4.510 3.525 4.850 5.280 ;
        RECT  1.670 3.820 2.015 5.280 ;
        RECT  0.180 3.870 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.025 ;
        RECT  0.170 1.795 1.815 2.025 ;
        RECT  0.780 1.795 1.815 2.135 ;
        RECT  0.780 1.795 1.120 3.085 ;
        RECT  2.045 1.175 2.940 1.515 ;
        RECT  0.260 3.235 0.600 3.575 ;
        RECT  2.045 1.175 2.275 3.575 ;
        RECT  0.260 3.345 3.450 3.575 ;
        RECT  3.110 3.345 3.450 3.665 ;
        RECT  6.695 1.240 7.035 1.845 ;
        RECT  5.345 1.615 7.035 1.845 ;
        RECT  5.345 1.615 5.625 2.095 ;
        RECT  5.345 1.615 5.605 2.120 ;
        RECT  6.725 1.240 7.035 2.540 ;
        RECT  6.725 2.310 8.125 2.540 ;
        RECT  7.785 2.310 8.125 2.650 ;
        RECT  6.560 2.540 6.955 2.880 ;
        RECT  2.790 2.500 3.130 3.115 ;
        RECT  6.560 2.540 6.790 3.295 ;
        RECT  2.790 2.885 4.425 3.115 ;
        RECT  4.195 3.065 6.790 3.295 ;
        RECT  6.235 0.780 7.495 1.010 ;
        RECT  4.885 1.070 5.245 1.385 ;
        RECT  6.235 0.780 6.465 1.385 ;
        RECT  4.885 1.155 6.465 1.385 ;
        RECT  4.885 1.070 5.240 1.410 ;
        RECT  7.265 0.780 7.495 1.870 ;
        RECT  7.265 1.640 8.565 1.870 ;
        RECT  2.505 1.745 3.675 1.975 ;
        RECT  8.225 1.750 8.690 1.980 ;
        RECT  2.505 1.745 2.790 2.085 ;
        RECT  3.445 1.745 3.675 2.655 ;
        RECT  3.445 2.290 3.900 2.655 ;
        RECT  3.445 2.425 5.115 2.655 ;
        RECT  4.885 1.070 5.115 2.655 ;
        RECT  8.460 1.750 8.690 3.080 ;
        RECT  4.905 2.550 5.350 2.835 ;
        RECT  8.460 2.740 8.800 3.080 ;
        RECT  8.505 1.070 9.225 1.410 ;
        RECT  8.995 1.070 9.225 2.460 ;
        RECT  9.035 2.635 10.830 2.975 ;
        RECT  9.035 2.230 9.265 3.550 ;
        RECT  8.380 3.320 9.265 3.550 ;
        RECT  8.380 3.320 8.720 4.250 ;
        RECT  9.455 1.180 11.080 1.410 ;
        RECT  9.455 1.180 9.795 1.720 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  11.070 1.695 11.570 2.500 ;
        RECT  11.070 2.160 11.725 2.500 ;
        RECT  11.070 1.695 11.300 3.435 ;
        RECT  9.970 3.205 11.300 3.435 ;
        RECT  9.970 3.205 10.310 3.605 ;
        RECT  0.260 3.345 2.70 3.575 ;
        RECT  4.195 3.065 5.70 3.295 ;
    END
END DFRSX1

MACRO DFRSX0
    CLASS CORE ;
    FOREIGN DFRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.645 2.715 11.215 3.240 ;
        RECT  10.985 0.630 11.215 3.240 ;
        RECT  10.070 0.630 11.215 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.760 2.220 4.285 2.685 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.360 2.210 9.955 2.630 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.502  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.445 1.170 11.845 3.765 ;
        END
    END QN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.630 2.135 6.175 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.645 3.515 10.985 5.280 ;
        RECT  8.690 3.635 9.030 5.280 ;
        RECT  6.095 3.630 6.435 5.280 ;
        RECT  5.050 3.910 5.390 5.280 ;
        RECT  4.120 3.910 4.460 5.280 ;
        RECT  1.470 3.360 1.810 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  11.450 -0.400 11.790 0.710 ;
        RECT  8.970 -0.400 9.315 0.970 ;
        RECT  7.140 -0.400 7.425 0.970 ;
        RECT  5.190 -0.400 5.475 0.970 ;
        RECT  3.890 -0.400 4.230 0.990 ;
        RECT  1.300 -0.400 1.640 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.270 0.630 0.610 1.930 ;
        RECT  0.115 1.700 1.905 1.930 ;
        RECT  1.620 1.700 1.905 2.080 ;
        RECT  0.115 1.700 0.345 3.060 ;
        RECT  0.115 2.770 1.080 3.060 ;
        RECT  0.740 2.770 1.080 3.700 ;
        RECT  2.690 1.165 3.030 1.505 ;
        RECT  2.135 1.210 3.030 1.505 ;
        RECT  0.575 2.200 0.860 2.540 ;
        RECT  2.135 1.210 2.365 2.540 ;
        RECT  0.575 2.310 2.365 2.540 ;
        RECT  2.040 2.310 2.270 4.140 ;
        RECT  2.040 3.910 3.120 4.140 ;
        RECT  2.780 3.910 3.120 4.250 ;
        RECT  6.165 1.270 6.450 1.905 ;
        RECT  4.975 2.160 5.315 2.500 ;
        RECT  6.405 1.675 6.635 3.200 ;
        RECT  5.085 2.860 7.385 3.200 ;
        RECT  2.500 2.840 2.840 3.675 ;
        RECT  5.085 2.160 5.315 3.675 ;
        RECT  2.500 3.445 5.315 3.675 ;
        RECT  5.705 0.810 6.910 1.040 ;
        RECT  6.680 0.810 6.910 1.445 ;
        RECT  5.705 0.810 5.935 1.610 ;
        RECT  4.515 1.270 5.935 1.610 ;
        RECT  2.595 1.735 4.745 1.965 ;
        RECT  2.595 1.735 3.510 2.080 ;
        RECT  6.865 1.215 7.095 2.460 ;
        RECT  6.865 2.120 8.000 2.460 ;
        RECT  4.515 1.270 4.745 3.200 ;
        RECT  3.170 1.735 3.510 3.180 ;
        RECT  4.450 2.860 4.790 3.200 ;
        RECT  7.715 2.120 8.000 3.425 ;
        RECT  7.940 0.630 8.460 0.970 ;
        RECT  8.230 2.880 9.955 3.110 ;
        RECT  9.640 2.880 9.955 3.220 ;
        RECT  8.230 0.630 8.460 3.970 ;
        RECT  7.435 3.655 8.460 3.970 ;
        RECT  8.690 1.690 10.410 1.920 ;
        RECT  10.070 1.310 10.410 1.920 ;
        RECT  8.690 1.690 9.030 2.105 ;
        RECT  10.185 1.830 10.755 2.170 ;
        RECT  10.185 1.830 10.415 3.970 ;
        RECT  9.510 3.630 10.415 3.970 ;
        RECT  5.085 2.860 6.60 3.200 ;
        RECT  2.500 3.445 4.50 3.675 ;
        RECT  2.595 1.735 3.80 1.965 ;
    END
END DFRSX0

MACRO DFRSQX4
    CLASS CORE ;
    FOREIGN DFRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.600 1.130 14.940 4.130 ;
        RECT  13.280 2.250 14.940 2.630 ;
        RECT  13.280 0.790 13.620 2.630 ;
        RECT  13.160 2.890 13.510 4.100 ;
        RECT  13.280 0.790 13.510 4.100 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.110 1.640 11.845 2.020 ;
        RECT  11.110 1.640 11.450 2.090 ;
        END
    END SN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.660 6.910 2.160 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  14.040 -0.400 14.380 0.720 ;
        RECT  12.520 -0.400 12.860 0.710 ;
        RECT  10.825 -0.400 11.165 0.910 ;
        RECT  8.060 -0.400 8.345 1.320 ;
        RECT  6.105 -0.400 6.445 0.970 ;
        RECT  1.580 -0.400 2.815 0.710 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  13.880 2.890 14.220 5.280 ;
        RECT  12.400 4.160 12.740 5.280 ;
        RECT  11.015 3.540 11.355 5.280 ;
        RECT  8.875 3.850 9.215 5.280 ;
        RECT  6.455 2.910 6.755 5.280 ;
        RECT  2.410 3.965 2.750 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 3.275 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.505 1.190 4.095 1.530 ;
        RECT  1.835 2.325 3.735 2.665 ;
        RECT  3.505 1.190 3.735 3.275 ;
        RECT  3.505 2.935 3.985 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.705 3.735 ;
        RECT  4.365 2.980 4.705 3.735 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  3.045 0.700 4.555 0.930 ;
        RECT  4.325 0.700 4.555 1.550 ;
        RECT  3.045 0.700 3.275 1.520 ;
        RECT  0.780 1.290 3.275 1.520 ;
        RECT  4.325 1.320 4.910 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.570 1.320 4.910 1.660 ;
        RECT  6.675 0.775 7.830 1.005 ;
        RECT  4.785 0.735 5.710 1.075 ;
        RECT  5.480 0.735 5.710 3.195 ;
        RECT  6.675 0.775 6.905 1.430 ;
        RECT  5.480 1.200 6.905 1.430 ;
        RECT  7.600 0.775 7.830 1.910 ;
        RECT  7.600 1.680 9.255 1.910 ;
        RECT  8.915 1.680 9.255 2.020 ;
        RECT  5.480 1.200 5.765 3.195 ;
        RECT  7.135 1.240 7.370 1.580 ;
        RECT  3.965 1.840 4.275 2.180 ;
        RECT  3.965 1.950 5.250 2.180 ;
        RECT  7.140 1.240 7.370 2.860 ;
        RECT  7.140 2.340 7.995 2.680 ;
        RECT  9.585 1.520 9.870 2.680 ;
        RECT  5.995 2.450 9.870 2.680 ;
        RECT  7.135 2.450 7.475 2.860 ;
        RECT  4.935 1.950 5.250 3.655 ;
        RECT  8.345 3.390 9.965 3.620 ;
        RECT  7.135 2.450 7.365 3.855 ;
        RECT  5.995 2.450 6.225 3.655 ;
        RECT  4.935 3.425 6.225 3.655 ;
        RECT  8.345 3.390 8.575 3.855 ;
        RECT  7.135 3.625 8.575 3.855 ;
        RECT  9.625 3.390 9.965 4.000 ;
        RECT  9.155 0.920 9.495 1.290 ;
        RECT  9.155 1.060 10.330 1.290 ;
        RECT  11.925 2.370 12.265 2.710 ;
        RECT  10.100 2.480 12.265 2.710 ;
        RECT  7.795 2.930 10.425 3.160 ;
        RECT  10.100 1.060 10.330 3.160 ;
        RECT  7.685 3.110 8.025 3.395 ;
        RECT  10.195 2.480 10.425 3.880 ;
        RECT  10.195 3.540 10.535 3.880 ;
        RECT  10.560 1.140 12.360 1.370 ;
        RECT  10.560 1.140 10.845 1.480 ;
        RECT  12.020 1.250 12.725 1.480 ;
        RECT  12.495 1.250 12.725 3.170 ;
        RECT  11.735 2.940 12.725 3.170 ;
        RECT  11.735 2.940 12.075 3.760 ;
        RECT  2.030 3.505 3.20 3.735 ;
        RECT  0.180 3.600 1.30 3.830 ;
        RECT  0.780 1.290 2.20 1.520 ;
        RECT  5.995 2.450 8.50 2.680 ;
        RECT  10.100 2.480 11.10 2.710 ;
        RECT  7.795 2.930 9.40 3.160 ;
    END
END DFRSQX4

MACRO DFRSQX2
    CLASS CORE ;
    FOREIGN DFRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.180 11.860 3.550 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.760 2.075 6.175 2.660 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.800 2.250 10.585 2.735 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 1.630 4.400 2.110 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  10.960 3.995 12.420 5.280 ;
        RECT  9.425 3.425 9.765 5.280 ;
        RECT  6.940 3.470 7.280 5.280 ;
        RECT  5.640 3.525 5.980 5.280 ;
        RECT  4.340 3.525 4.680 5.280 ;
        RECT  1.700 3.910 2.550 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.960 -0.400 12.420 0.720 ;
        RECT  9.205 -0.400 9.545 1.090 ;
        RECT  7.280 -0.400 7.620 0.890 ;
        RECT  5.270 -0.400 5.610 0.925 ;
        RECT  3.640 -0.400 3.980 0.725 ;
        RECT  1.130 -0.400 1.470 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.700 ;
        RECT  0.115 2.585 2.040 2.815 ;
        RECT  1.730 2.585 2.040 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  1.700 1.035 2.780 1.325 ;
        RECT  1.700 1.035 1.930 2.355 ;
        RECT  1.700 2.125 2.500 2.355 ;
        RECT  0.575 3.100 0.915 3.440 ;
        RECT  2.270 2.125 2.500 3.575 ;
        RECT  0.575 3.210 2.500 3.440 ;
        RECT  2.270 3.345 3.350 3.575 ;
        RECT  3.010 3.345 3.350 3.685 ;
        RECT  6.300 1.240 6.590 1.845 ;
        RECT  5.090 1.615 6.635 1.845 ;
        RECT  5.090 1.615 5.430 2.100 ;
        RECT  6.405 1.615 6.635 3.295 ;
        RECT  6.405 2.280 8.035 2.510 ;
        RECT  7.695 2.280 8.035 2.605 ;
        RECT  2.730 2.310 3.060 2.650 ;
        RECT  2.830 2.310 3.060 3.115 ;
        RECT  6.400 2.780 6.740 3.295 ;
        RECT  2.830 2.885 4.330 3.115 ;
        RECT  6.405 2.280 6.740 3.295 ;
        RECT  4.100 3.065 6.740 3.295 ;
        RECT  5.840 0.780 7.050 1.010 ;
        RECT  6.820 0.780 7.050 1.390 ;
        RECT  5.840 0.780 6.070 1.385 ;
        RECT  4.510 1.155 6.070 1.385 ;
        RECT  6.820 1.160 7.435 1.390 ;
        RECT  4.510 1.070 4.850 1.410 ;
        RECT  2.160 1.555 2.500 1.895 ;
        RECT  7.205 1.160 7.435 2.010 ;
        RECT  7.205 1.670 7.545 2.010 ;
        RECT  2.160 1.665 3.620 1.895 ;
        RECT  7.205 1.780 8.495 2.010 ;
        RECT  3.390 1.665 3.620 2.655 ;
        RECT  3.390 2.290 3.730 2.655 ;
        RECT  4.630 1.155 4.860 2.835 ;
        RECT  3.390 2.425 4.860 2.655 ;
        RECT  4.630 2.550 5.220 2.835 ;
        RECT  8.265 1.780 8.495 3.065 ;
        RECT  7.635 2.835 8.495 3.065 ;
        RECT  7.635 2.835 7.865 4.040 ;
        RECT  7.635 3.810 8.795 4.040 ;
        RECT  8.455 3.810 8.795 4.100 ;
        RECT  8.175 0.630 8.955 0.950 ;
        RECT  8.725 2.965 10.775 3.195 ;
        RECT  10.435 2.965 10.775 3.305 ;
        RECT  8.725 0.630 8.955 3.580 ;
        RECT  8.095 3.295 8.955 3.580 ;
        RECT  10.235 0.680 10.575 2.020 ;
        RECT  9.185 1.790 11.235 2.020 ;
        RECT  9.185 1.790 9.470 2.700 ;
        RECT  11.005 1.790 11.235 3.765 ;
        RECT  10.200 3.535 11.235 3.765 ;
        RECT  10.200 3.535 10.540 4.070 ;
        RECT  4.100 3.065 5.80 3.295 ;
        RECT  8.725 2.965 9.40 3.195 ;
        RECT  9.185 1.790 10.40 2.020 ;
    END
END DFRSQX2

MACRO DFRSQX1
    CLASS CORE ;
    FOREIGN DFRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.230 1.640 4.570 2.085 ;
        RECT  3.905 1.640 4.570 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.955 2.075 6.415 2.360 ;
        RECT  5.795 2.250 6.175 2.630 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.640 10.585 2.305 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.530 2.400 12.475 2.630 ;
        RECT  12.095 2.250 12.475 2.630 ;
        RECT  12.095 1.235 12.325 2.630 ;
        RECT  11.380 1.235 12.325 1.465 ;
        RECT  11.270 3.665 11.760 4.005 ;
        RECT  11.530 2.400 11.760 4.005 ;
        RECT  11.380 0.700 11.610 1.465 ;
        RECT  11.270 0.700 11.610 1.040 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.990 -0.400 12.330 1.005 ;
        RECT  10.015 -0.400 10.355 0.880 ;
        RECT  7.725 -0.400 8.065 0.790 ;
        RECT  5.665 -0.400 6.005 0.925 ;
        RECT  4.165 -0.400 4.505 1.410 ;
        RECT  1.340 -0.400 1.680 1.565 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.990 3.330 12.330 5.280 ;
        RECT  10.570 4.005 10.910 5.280 ;
        RECT  9.210 3.910 9.550 5.280 ;
        RECT  7.110 3.320 7.450 5.280 ;
        RECT  5.810 3.525 6.150 5.280 ;
        RECT  4.510 3.525 4.850 5.280 ;
        RECT  1.670 3.820 2.015 5.280 ;
        RECT  0.180 3.870 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.025 ;
        RECT  0.170 1.795 1.815 2.025 ;
        RECT  1.475 1.795 1.815 2.135 ;
        RECT  0.780 1.795 1.120 3.085 ;
        RECT  2.045 1.175 2.940 1.515 ;
        RECT  0.260 3.235 0.600 3.575 ;
        RECT  2.045 1.175 2.275 3.575 ;
        RECT  0.260 3.345 3.450 3.575 ;
        RECT  3.110 3.345 3.450 3.665 ;
        RECT  6.695 1.240 7.035 1.580 ;
        RECT  6.695 1.240 6.955 1.845 ;
        RECT  5.345 1.615 6.955 1.845 ;
        RECT  5.345 1.615 5.625 2.095 ;
        RECT  5.345 1.615 5.605 2.120 ;
        RECT  6.725 2.310 8.125 2.540 ;
        RECT  7.785 2.310 8.125 2.650 ;
        RECT  6.725 1.240 6.955 2.880 ;
        RECT  2.790 2.500 3.130 3.115 ;
        RECT  6.560 2.540 6.790 3.295 ;
        RECT  2.790 2.885 4.425 3.115 ;
        RECT  4.195 3.065 6.790 3.295 ;
        RECT  6.235 0.780 7.495 1.010 ;
        RECT  4.885 1.070 5.245 1.385 ;
        RECT  6.235 0.780 6.465 1.385 ;
        RECT  4.885 1.155 6.465 1.385 ;
        RECT  4.885 1.070 5.240 1.410 ;
        RECT  7.265 0.780 7.495 1.870 ;
        RECT  7.265 1.640 8.565 1.870 ;
        RECT  8.225 1.750 8.690 1.980 ;
        RECT  2.505 1.745 3.675 2.085 ;
        RECT  3.445 1.745 3.675 2.655 ;
        RECT  3.445 2.290 3.900 2.655 ;
        RECT  3.445 2.425 5.115 2.655 ;
        RECT  4.885 1.070 5.115 2.655 ;
        RECT  8.460 1.750 8.690 3.080 ;
        RECT  4.905 2.550 5.350 2.835 ;
        RECT  8.460 2.740 8.800 3.080 ;
        RECT  8.505 1.070 9.225 1.410 ;
        RECT  8.995 1.070 9.225 2.460 ;
        RECT  9.035 2.635 10.830 2.865 ;
        RECT  10.490 2.635 10.830 2.975 ;
        RECT  9.035 2.230 9.265 3.550 ;
        RECT  8.380 3.320 9.265 3.550 ;
        RECT  8.380 3.320 8.720 4.250 ;
        RECT  9.455 1.180 11.080 1.410 ;
        RECT  9.455 1.180 9.795 1.720 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  11.070 1.695 11.570 1.980 ;
        RECT  11.070 1.695 11.300 3.435 ;
        RECT  9.970 3.205 11.300 3.435 ;
        RECT  9.970 3.205 10.310 3.605 ;
        RECT  0.260 3.345 2.30 3.575 ;
        RECT  4.195 3.065 5.20 3.295 ;
    END
END DFRSQX1

MACRO DFRSQX0
    CLASS CORE ;
    FOREIGN DFRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.542  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.670 2.715 11.215 3.240 ;
        RECT  10.985 0.630 11.215 3.240 ;
        RECT  10.200 0.630 11.215 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.760 2.220 4.285 2.685 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.360 2.210 9.955 2.630 ;
        END
    END SN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.630 2.135 6.175 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.670 3.515 11.010 5.280 ;
        RECT  8.690 3.635 9.030 5.280 ;
        RECT  6.095 3.630 6.435 5.280 ;
        RECT  5.050 3.910 5.390 5.280 ;
        RECT  4.120 3.910 4.460 5.280 ;
        RECT  1.470 3.360 1.810 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  8.970 -0.400 9.310 1.420 ;
        RECT  7.140 -0.400 7.425 0.970 ;
        RECT  5.190 -0.400 5.475 0.970 ;
        RECT  3.890 -0.400 4.230 0.990 ;
        RECT  1.300 -0.400 1.640 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.270 0.630 0.610 1.930 ;
        RECT  0.115 1.700 1.905 1.930 ;
        RECT  1.620 1.700 1.905 2.080 ;
        RECT  0.115 1.700 0.345 3.060 ;
        RECT  0.115 2.770 1.080 3.060 ;
        RECT  0.740 2.770 1.080 3.700 ;
        RECT  2.690 1.165 3.030 1.505 ;
        RECT  2.135 1.275 3.030 1.505 ;
        RECT  0.575 2.200 0.860 2.540 ;
        RECT  2.135 1.275 2.365 2.540 ;
        RECT  0.575 2.310 2.365 2.540 ;
        RECT  2.040 2.310 2.270 4.140 ;
        RECT  2.040 3.910 3.120 4.140 ;
        RECT  2.780 3.910 3.120 4.250 ;
        RECT  6.165 1.270 6.450 1.905 ;
        RECT  4.975 2.160 5.315 2.500 ;
        RECT  6.405 1.675 6.635 3.200 ;
        RECT  2.500 2.840 2.840 3.180 ;
        RECT  5.085 2.860 7.385 3.200 ;
        RECT  2.610 2.840 2.840 3.675 ;
        RECT  5.085 2.160 5.315 3.675 ;
        RECT  2.610 3.445 5.315 3.675 ;
        RECT  5.705 0.810 6.910 1.040 ;
        RECT  6.680 0.810 6.910 1.445 ;
        RECT  5.705 0.810 5.935 1.610 ;
        RECT  4.515 1.270 5.935 1.610 ;
        RECT  2.595 1.735 4.745 1.965 ;
        RECT  2.595 1.735 3.510 2.080 ;
        RECT  6.865 1.215 7.095 2.460 ;
        RECT  6.865 2.120 8.000 2.460 ;
        RECT  4.515 1.270 4.745 3.200 ;
        RECT  3.170 1.735 3.510 3.180 ;
        RECT  4.450 2.860 4.790 3.200 ;
        RECT  7.715 2.120 8.000 3.425 ;
        RECT  7.940 0.630 8.460 0.970 ;
        RECT  8.230 2.880 9.980 3.110 ;
        RECT  9.640 2.880 9.980 3.220 ;
        RECT  8.230 0.630 8.460 3.970 ;
        RECT  7.435 3.655 8.460 3.970 ;
        RECT  10.200 1.310 10.540 1.650 ;
        RECT  10.200 1.310 10.440 1.920 ;
        RECT  8.690 1.690 10.440 1.920 ;
        RECT  8.690 1.690 9.030 2.105 ;
        RECT  10.210 1.310 10.440 3.970 ;
        RECT  9.510 3.630 10.440 3.970 ;
        RECT  5.085 2.860 6.50 3.200 ;
        RECT  2.610 3.445 4.00 3.675 ;
        RECT  2.595 1.735 3.40 1.965 ;
    END
END DFRSQX0

MACRO DFRRX4
    CLASS CORE ;
    FOREIGN DFRRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.002  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.380 1.130 18.775 3.175 ;
        RECT  17.180 2.250 18.775 2.630 ;
        RECT  17.180 2.250 17.560 3.195 ;
        RECT  17.180 1.130 17.410 3.195 ;
        RECT  16.940 1.130 17.410 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.078  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.880 16.950 3.220 ;
        RECT  16.720 1.700 16.950 3.220 ;
        RECT  14.170 1.700 16.950 1.930 ;
        RECT  15.500 1.130 15.840 1.930 ;
        RECT  14.615 2.640 14.995 4.180 ;
        RECT  14.170 1.130 14.400 1.930 ;
        RECT  14.060 1.130 14.400 1.470 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.290 1.640 13.105 2.020 ;
        RECT  12.290 1.640 12.630 2.190 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.660 7.850 2.225 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.760 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  17.660 -0.400 18.000 1.470 ;
        RECT  16.220 -0.400 16.560 1.470 ;
        RECT  14.780 -0.400 15.120 1.470 ;
        RECT  12.800 -0.400 13.140 0.710 ;
        RECT  7.230 -0.400 7.515 0.970 ;
        RECT  1.750 -0.400 3.225 0.655 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  17.800 3.510 18.140 5.280 ;
        RECT  16.640 3.580 16.980 5.280 ;
        RECT  15.390 3.870 15.730 5.280 ;
        RECT  13.870 4.110 14.210 5.280 ;
        RECT  11.490 3.760 12.950 5.280 ;
        RECT  9.315 4.170 9.655 5.280 ;
        RECT  6.825 3.925 7.165 5.280 ;
        RECT  2.410 3.985 3.245 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.805 1.920 2.090 ;
        RECT  1.375 1.860 3.420 2.090 ;
        RECT  3.190 1.860 3.420 2.800 ;
        RECT  3.190 2.460 3.530 2.800 ;
        RECT  1.375 1.805 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.780 1.345 3.935 1.575 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  2.325 1.345 3.935 1.630 ;
        RECT  3.645 1.345 3.935 1.695 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.525 5.200 3.755 ;
        RECT  4.860 3.010 5.200 3.755 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  4.165 1.160 5.210 1.500 ;
        RECT  1.835 2.325 2.580 2.665 ;
        RECT  4.165 1.160 4.395 3.295 ;
        RECT  2.240 2.325 2.580 3.295 ;
        RECT  4.140 2.955 4.480 3.295 ;
        RECT  2.240 3.065 4.480 3.295 ;
        RECT  0.180 0.640 0.520 1.015 ;
        RECT  3.520 0.700 5.670 0.930 ;
        RECT  0.180 0.785 1.520 1.015 ;
        RECT  1.290 0.885 3.750 1.115 ;
        RECT  5.440 0.700 5.670 1.640 ;
        RECT  5.440 1.320 6.025 1.640 ;
        RECT  7.745 0.775 8.895 1.005 ;
        RECT  5.900 0.735 6.770 1.090 ;
        RECT  6.255 0.735 6.770 1.430 ;
        RECT  7.745 0.775 7.975 1.430 ;
        RECT  6.255 1.200 7.975 1.430 ;
        RECT  8.665 0.775 8.895 2.090 ;
        RECT  8.665 1.860 10.330 2.090 ;
        RECT  9.990 1.860 10.330 2.200 ;
        RECT  6.255 0.735 6.485 3.235 ;
        RECT  6.050 2.895 6.485 3.235 ;
        RECT  4.625 1.820 4.935 2.175 ;
        RECT  4.625 1.890 5.810 2.175 ;
        RECT  8.205 1.240 8.435 2.805 ;
        RECT  8.205 2.340 8.685 2.805 ;
        RECT  8.205 2.520 11.000 2.805 ;
        RECT  10.660 1.670 11.000 2.805 ;
        RECT  7.585 2.575 11.000 2.805 ;
        RECT  7.585 2.575 7.925 2.915 ;
        RECT  5.470 1.890 5.810 3.695 ;
        RECT  5.470 3.465 7.815 3.695 ;
        RECT  7.585 2.575 7.815 3.940 ;
        RECT  7.585 3.710 10.170 3.940 ;
        RECT  9.940 3.710 10.170 4.250 ;
        RECT  9.940 3.965 10.280 4.250 ;
        RECT  9.125 0.630 12.340 0.860 ;
        RECT  11.530 0.630 12.340 0.950 ;
        RECT  9.125 0.630 9.420 1.500 ;
        RECT  10.230 1.100 10.570 1.440 ;
        RECT  10.230 1.210 11.460 1.440 ;
        RECT  13.140 2.310 13.480 2.650 ;
        RECT  11.230 2.420 13.480 2.650 ;
        RECT  12.050 2.420 12.390 3.150 ;
        RECT  11.230 1.210 11.460 3.395 ;
        RECT  8.125 3.165 11.460 3.395 ;
        RECT  8.125 3.165 8.465 3.480 ;
        RECT  10.485 3.165 10.800 3.860 ;
        RECT  10.510 3.165 10.800 3.890 ;
        RECT  11.690 1.180 13.700 1.410 ;
        RECT  13.360 1.110 13.700 1.905 ;
        RECT  11.690 1.180 11.975 1.730 ;
        RECT  13.360 1.675 13.940 1.905 ;
        RECT  13.710 2.180 16.480 2.410 ;
        RECT  16.140 2.180 16.480 2.650 ;
        RECT  13.710 1.675 13.940 3.110 ;
        RECT  13.310 2.880 13.940 3.110 ;
        RECT  13.310 2.880 13.650 3.700 ;
        RECT  1.375 1.860 2.80 2.090 ;
        RECT  0.780 1.345 2.40 1.575 ;
        RECT  2.030 3.525 4.90 3.755 ;
        RECT  0.180 3.600 1.40 3.830 ;
        RECT  2.240 3.065 3.90 3.295 ;
        RECT  3.520 0.700 4.30 0.930 ;
        RECT  1.290 0.885 2.20 1.115 ;
        RECT  8.205 2.520 10.80 2.805 ;
        RECT  7.585 2.575 10.60 2.805 ;
        RECT  5.470 3.465 6.30 3.695 ;
        RECT  7.585 3.710 9.20 3.940 ;
        RECT  9.125 0.630 11.50 0.860 ;
        RECT  11.230 2.420 12.00 2.650 ;
        RECT  8.125 3.165 10.40 3.395 ;
        RECT  11.690 1.180 12.60 1.410 ;
        RECT  13.710 2.180 15.50 2.410 ;
    END
END DFRRX4

MACRO DFRRX2
    CLASS CORE ;
    FOREIGN DFRRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 1.240 13.750 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.090 2.860 13.105 3.090 ;
        RECT  12.875 0.950 13.105 3.090 ;
        RECT  12.090 0.950 13.105 1.180 ;
        RECT  12.090 2.860 12.475 4.180 ;
        RECT  12.090 0.820 12.430 1.180 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.080 1.940 10.585 2.630 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.075 6.390 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.400 1.640 4.915 2.120 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  12.850 3.950 14.310 5.280 ;
        RECT  11.370 3.785 11.710 5.280 ;
        RECT  9.620 3.860 9.960 5.280 ;
        RECT  7.200 3.660 7.540 5.280 ;
        RECT  5.900 3.525 6.240 5.280 ;
        RECT  4.600 3.525 4.940 5.280 ;
        RECT  1.470 3.805 2.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  12.850 -0.400 14.310 0.720 ;
        RECT  11.330 -0.400 11.670 0.720 ;
        RECT  10.430 -0.400 10.770 0.710 ;
        RECT  5.390 -0.400 5.730 0.925 ;
        RECT  0.780 -0.400 1.120 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.360 0.520 2.510 ;
        RECT  0.115 2.280 1.905 2.510 ;
        RECT  1.620 2.280 1.905 2.620 ;
        RECT  0.115 2.280 0.345 4.070 ;
        RECT  0.115 3.730 0.620 4.070 ;
        RECT  2.700 1.305 3.040 1.645 ;
        RECT  2.135 1.415 3.040 1.645 ;
        RECT  0.575 2.850 2.365 3.190 ;
        RECT  2.135 1.415 2.365 3.575 ;
        RECT  2.135 3.345 3.630 3.575 ;
        RECT  3.290 3.345 3.630 3.685 ;
        RECT  1.580 0.630 4.240 0.950 ;
        RECT  1.580 0.630 1.920 1.090 ;
        RECT  6.420 1.240 6.710 1.845 ;
        RECT  5.145 1.615 6.850 1.845 ;
        RECT  5.145 1.615 5.450 2.195 ;
        RECT  6.620 1.615 6.850 3.295 ;
        RECT  7.920 2.360 8.260 2.700 ;
        RECT  6.620 2.470 8.260 2.700 ;
        RECT  3.010 2.505 3.350 3.115 ;
        RECT  3.010 2.885 4.910 3.115 ;
        RECT  6.620 2.470 7.000 3.295 ;
        RECT  4.680 3.065 7.000 3.295 ;
        RECT  5.960 0.780 7.310 1.010 ;
        RECT  4.630 1.155 6.190 1.385 ;
        RECT  5.960 0.780 6.190 1.385 ;
        RECT  4.630 1.070 4.970 1.410 ;
        RECT  3.680 1.180 4.970 1.410 ;
        RECT  7.080 0.780 7.310 1.980 ;
        RECT  7.080 1.750 7.660 1.980 ;
        RECT  7.320 1.860 8.740 2.090 ;
        RECT  2.595 1.880 3.910 2.220 ;
        RECT  3.680 1.180 3.910 2.655 ;
        RECT  3.680 2.315 4.020 2.655 ;
        RECT  3.680 2.425 5.480 2.655 ;
        RECT  8.510 1.860 8.740 3.130 ;
        RECT  5.140 2.425 5.480 2.835 ;
        RECT  8.510 2.790 9.010 3.130 ;
        RECT  7.540 0.630 10.010 0.970 ;
        RECT  9.670 0.630 10.010 1.040 ;
        RECT  8.440 1.210 9.200 1.550 ;
        RECT  8.970 1.210 9.200 2.200 ;
        RECT  8.970 1.970 9.550 2.200 ;
        RECT  9.320 2.860 11.135 3.090 ;
        RECT  10.795 2.750 11.135 3.095 ;
        RECT  10.180 2.860 11.135 3.095 ;
        RECT  10.180 2.860 10.520 3.200 ;
        RECT  9.320 1.970 9.550 3.630 ;
        RECT  8.385 3.400 9.550 3.630 ;
        RECT  8.385 3.400 8.725 3.825 ;
        RECT  9.430 1.400 11.670 1.630 ;
        RECT  9.430 1.400 9.770 1.740 ;
        RECT  11.330 1.400 11.670 1.980 ;
        RECT  11.440 2.120 12.645 2.460 ;
        RECT  11.440 1.400 11.670 3.555 ;
        RECT  10.760 3.325 11.670 3.555 ;
        RECT  10.760 3.325 10.990 4.125 ;
        RECT  10.650 3.785 10.990 4.125 ;
        RECT  1.580 0.630 3.10 0.950 ;
        RECT  4.680 3.065 6.40 3.295 ;
        RECT  7.540 0.630 9.60 0.970 ;
        RECT  9.430 1.400 10.40 1.630 ;
    END
END DFRRX2

MACRO DFRRX1
    CLASS CORE ;
    FOREIGN DFRRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.655 2.025 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.955 2.075 6.490 2.360 ;
        RECT  5.795 2.250 6.175 2.630 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.050 1.640 10.610 2.085 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.678  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 2.250 12.475 2.630 ;
        RECT  11.530 2.870 12.325 3.100 ;
        RECT  12.095 1.235 12.325 3.100 ;
        RECT  11.380 1.235 12.325 1.465 ;
        RECT  11.270 3.435 11.760 3.720 ;
        RECT  11.530 2.870 11.760 3.720 ;
        RECT  11.380 0.700 11.610 1.465 ;
        RECT  11.270 0.700 11.610 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 0.820 13.105 4.180 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.990 -0.400 12.330 1.005 ;
        RECT  10.470 -0.400 10.810 0.950 ;
        RECT  5.725 -0.400 6.065 0.925 ;
        RECT  0.915 -0.400 1.255 1.395 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  11.990 3.330 12.330 5.280 ;
        RECT  9.800 3.840 10.140 5.280 ;
        RECT  7.185 3.480 7.525 5.280 ;
        RECT  5.885 3.525 6.225 5.280 ;
        RECT  4.585 3.525 4.925 5.280 ;
        RECT  1.940 3.840 2.280 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.215 0.645 0.555 2.350 ;
        RECT  0.115 2.120 1.950 2.350 ;
        RECT  1.665 2.120 1.950 2.460 ;
        RECT  0.115 2.120 0.345 3.790 ;
        RECT  0.115 3.450 0.760 3.790 ;
        RECT  2.180 1.090 3.205 1.325 ;
        RECT  0.575 2.855 1.555 3.195 ;
        RECT  1.220 2.855 1.555 4.180 ;
        RECT  2.180 1.090 2.410 3.575 ;
        RECT  1.220 3.345 3.525 3.575 ;
        RECT  3.185 3.345 3.525 3.665 ;
        RECT  1.220 3.345 1.560 4.180 ;
        RECT  1.635 0.630 4.605 0.860 ;
        RECT  4.265 0.630 4.605 1.410 ;
        RECT  1.635 0.630 1.950 1.450 ;
        RECT  5.345 1.615 7.040 1.845 ;
        RECT  5.345 1.615 5.625 2.095 ;
        RECT  5.345 1.615 5.605 2.120 ;
        RECT  6.755 1.240 7.040 2.690 ;
        RECT  6.755 2.460 8.200 2.690 ;
        RECT  7.860 2.460 8.200 2.800 ;
        RECT  2.905 2.500 3.215 3.115 ;
        RECT  6.635 2.720 6.985 3.295 ;
        RECT  2.905 2.885 4.490 3.115 ;
        RECT  6.755 1.240 6.985 3.295 ;
        RECT  4.260 3.065 6.985 3.295 ;
        RECT  6.295 0.780 7.500 1.010 ;
        RECT  4.885 1.070 5.305 1.385 ;
        RECT  6.295 0.780 6.525 1.385 ;
        RECT  4.885 1.155 6.525 1.385 ;
        RECT  4.885 1.070 5.295 1.390 ;
        RECT  2.640 1.555 3.675 1.785 ;
        RECT  7.270 0.780 7.500 2.020 ;
        RECT  2.640 1.555 2.925 1.895 ;
        RECT  7.270 1.790 8.660 2.020 ;
        RECT  7.990 1.790 8.660 2.130 ;
        RECT  3.445 1.555 3.675 2.655 ;
        RECT  3.445 2.290 3.975 2.655 ;
        RECT  3.445 2.425 5.115 2.655 ;
        RECT  4.885 1.070 5.115 2.655 ;
        RECT  4.905 2.550 5.425 2.835 ;
        RECT  8.430 1.790 8.660 3.240 ;
        RECT  8.430 2.900 8.960 3.240 ;
        RECT  7.730 0.630 10.010 0.860 ;
        RECT  9.670 0.630 10.010 0.950 ;
        RECT  7.730 0.630 8.070 0.970 ;
        RECT  8.440 1.220 9.155 1.560 ;
        RECT  8.925 1.220 9.155 2.635 ;
        RECT  8.925 2.405 10.830 2.635 ;
        RECT  10.130 2.405 10.830 2.745 ;
        RECT  10.130 2.405 10.470 3.375 ;
        RECT  9.290 2.405 9.520 3.820 ;
        RECT  8.340 3.480 9.520 3.820 ;
        RECT  9.390 1.180 11.080 1.410 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  9.390 1.180 9.730 2.010 ;
        RECT  11.070 1.695 11.765 2.545 ;
        RECT  11.070 2.205 11.865 2.545 ;
        RECT  11.070 1.695 11.300 3.205 ;
        RECT  10.770 2.975 11.300 3.205 ;
        RECT  10.770 2.975 11.000 4.180 ;
        RECT  10.600 3.840 11.000 4.180 ;
        RECT  1.220 3.345 2.80 3.575 ;
        RECT  1.635 0.630 3.40 0.860 ;
        RECT  4.260 3.065 5.40 3.295 ;
        RECT  7.730 0.630 9.30 0.860 ;
    END
END DFRRX1

MACRO DFRRX0
    CLASS CORE ;
    FOREIGN DFRRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.577  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.315 2.860 11.875 3.350 ;
        RECT  11.645 0.630 11.875 3.350 ;
        RECT  11.180 0.630 11.875 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.245 4.550 2.630 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.500 2.250 10.025 2.815 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.441  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.105 1.170 12.475 4.150 ;
        END
    END QN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.200 6.365 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.315 3.810 11.655 5.280 ;
        RECT  9.245 3.910 9.580 5.280 ;
        RECT  6.650 3.630 6.990 5.280 ;
        RECT  4.490 3.910 5.765 5.280 ;
        RECT  0.980 3.520 1.920 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.105 -0.400 12.420 0.710 ;
        RECT  10.380 -0.400 10.720 0.950 ;
        RECT  5.710 -0.400 5.995 1.400 ;
        RECT  0.780 -0.400 1.120 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.970 ;
        RECT  0.115 1.740 2.015 1.970 ;
        RECT  1.730 1.740 2.015 2.460 ;
        RECT  0.115 1.360 0.345 3.860 ;
        RECT  0.115 3.520 0.520 3.860 ;
        RECT  2.245 1.285 3.150 1.590 ;
        RECT  0.630 2.200 0.970 3.060 ;
        RECT  0.630 2.720 2.475 3.060 ;
        RECT  2.245 1.285 2.475 4.140 ;
        RECT  2.245 3.910 3.490 4.140 ;
        RECT  3.110 3.910 3.490 4.250 ;
        RECT  1.580 0.825 4.550 1.055 ;
        RECT  1.580 0.825 1.920 1.510 ;
        RECT  4.210 0.825 4.550 1.545 ;
        RECT  5.285 2.160 5.565 2.500 ;
        RECT  6.685 1.230 6.945 3.200 ;
        RECT  2.870 2.840 3.210 3.180 ;
        RECT  5.335 2.860 7.940 3.200 ;
        RECT  2.920 2.840 3.210 3.675 ;
        RECT  5.335 2.160 5.565 3.675 ;
        RECT  2.920 3.445 5.565 3.675 ;
        RECT  6.225 0.765 7.405 0.995 ;
        RECT  4.825 1.230 5.250 1.905 ;
        RECT  4.825 1.675 6.455 1.905 ;
        RECT  6.225 0.765 6.455 1.905 ;
        RECT  3.445 1.775 5.055 2.005 ;
        RECT  7.175 0.765 7.405 2.530 ;
        RECT  2.705 1.835 3.675 2.180 ;
        RECT  7.175 2.170 8.555 2.530 ;
        RECT  3.445 1.775 3.675 3.180 ;
        RECT  4.825 1.230 5.055 3.200 ;
        RECT  3.445 2.860 3.880 3.180 ;
        RECT  4.765 2.860 5.105 3.200 ;
        RECT  8.270 2.170 8.555 3.450 ;
        RECT  7.635 0.630 9.850 0.860 ;
        RECT  7.635 0.630 7.920 0.970 ;
        RECT  9.510 0.630 9.850 0.970 ;
        RECT  8.480 1.170 8.820 1.510 ;
        RECT  8.785 3.125 10.625 3.465 ;
        RECT  8.785 1.280 9.015 3.970 ;
        RECT  7.950 3.680 9.015 3.970 ;
        RECT  9.430 1.690 11.415 1.920 ;
        RECT  9.430 1.690 9.770 2.020 ;
        RECT  11.065 1.360 11.415 2.220 ;
        RECT  10.855 1.690 11.085 4.155 ;
        RECT  10.065 3.925 11.085 4.155 ;
        RECT  10.065 3.925 10.405 4.250 ;
        RECT  1.580 0.825 3.20 1.055 ;
        RECT  5.335 2.860 6.80 3.200 ;
        RECT  2.920 3.445 4.80 3.675 ;
        RECT  7.635 0.630 8.80 0.860 ;
    END
END DFRRX0

MACRO DFRRSX4
    CLASS CORE ;
    FOREIGN DFRRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.105  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 1.130 19.980 3.295 ;
        RECT  18.345 2.250 19.980 2.630 ;
        RECT  18.345 2.250 18.685 3.295 ;
        RECT  18.345 1.130 18.575 3.295 ;
        RECT  18.200 1.130 18.575 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.135  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.635 3.010 18.065 3.240 ;
        RECT  17.835 1.700 18.065 3.240 ;
        RECT  15.580 1.700 18.065 1.930 ;
        RECT  17.075 3.010 17.415 3.350 ;
        RECT  16.760 1.130 17.100 1.930 ;
        RECT  15.635 2.860 16.255 3.240 ;
        RECT  15.635 2.860 15.975 4.030 ;
        RECT  15.580 1.130 15.810 1.930 ;
        RECT  15.320 1.130 15.810 1.470 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.905 1.640 14.365 2.525 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.250 13.485 2.630 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.660 8.495 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.470 ;
        RECT  17.480 -0.400 17.820 1.470 ;
        RECT  16.040 -0.400 16.380 1.470 ;
        RECT  13.430 -0.400 13.770 0.950 ;
        RECT  7.830 -0.400 8.115 0.970 ;
        RECT  2.255 -0.400 3.825 0.665 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  19.000 3.530 19.340 5.280 ;
        RECT  17.705 3.685 18.045 5.280 ;
        RECT  16.355 3.470 16.695 5.280 ;
        RECT  14.875 4.060 15.215 5.280 ;
        RECT  12.435 3.910 13.895 5.280 ;
        RECT  10.135 3.965 10.475 5.280 ;
        RECT  7.715 2.910 8.015 5.280 ;
        RECT  2.410 3.965 3.845 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.765 1.815 2.105 2.095 ;
        RECT  1.375 1.860 4.020 2.095 ;
        RECT  3.790 1.860 4.020 2.800 ;
        RECT  3.790 2.460 4.130 2.800 ;
        RECT  1.375 1.860 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.965 1.355 4.535 1.585 ;
        RECT  0.965 1.290 1.305 1.630 ;
        RECT  2.925 1.355 4.535 1.630 ;
        RECT  4.245 1.355 4.535 1.695 ;
        RECT  4.765 1.160 5.810 1.500 ;
        RECT  1.835 2.325 2.120 2.665 ;
        RECT  1.835 2.435 3.070 2.665 ;
        RECT  2.840 2.435 3.070 3.275 ;
        RECT  2.840 2.935 3.180 3.275 ;
        RECT  4.765 1.160 4.995 3.540 ;
        RECT  2.840 3.045 4.995 3.275 ;
        RECT  4.735 3.200 5.080 3.540 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.415 3.735 ;
        RECT  4.185 3.505 4.415 4.000 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  5.500 2.980 5.840 4.000 ;
        RECT  4.185 3.770 5.840 4.000 ;
        RECT  0.365 0.640 0.705 1.015 ;
        RECT  4.120 0.630 6.270 0.860 ;
        RECT  0.365 0.785 2.025 1.015 ;
        RECT  4.120 0.630 4.350 1.125 ;
        RECT  1.795 0.895 4.350 1.125 ;
        RECT  6.040 0.630 6.270 1.660 ;
        RECT  6.040 1.320 6.625 1.660 ;
        RECT  8.345 0.775 9.495 1.005 ;
        RECT  6.500 0.735 7.370 1.090 ;
        RECT  8.345 0.775 8.575 1.430 ;
        RECT  7.140 1.200 8.575 1.430 ;
        RECT  9.265 0.775 9.495 2.090 ;
        RECT  9.265 1.860 10.930 2.090 ;
        RECT  7.140 0.735 7.370 2.150 ;
        RECT  6.740 1.920 7.370 2.150 ;
        RECT  10.590 1.860 10.930 2.200 ;
        RECT  6.740 1.920 7.025 3.195 ;
        RECT  5.225 1.820 5.535 2.175 ;
        RECT  11.260 1.670 11.600 2.010 ;
        RECT  5.225 1.945 6.510 2.175 ;
        RECT  8.805 1.240 9.035 2.680 ;
        RECT  8.805 2.340 9.505 2.680 ;
        RECT  11.260 1.670 11.490 2.680 ;
        RECT  7.255 2.450 11.490 2.680 ;
        RECT  8.395 2.450 8.735 2.860 ;
        RECT  6.170 1.945 6.510 3.655 ;
        RECT  8.395 2.450 8.625 3.855 ;
        RECT  7.255 2.450 7.485 3.655 ;
        RECT  6.170 3.425 7.485 3.655 ;
        RECT  9.605 3.505 11.225 3.735 ;
        RECT  8.395 3.625 9.835 3.855 ;
        RECT  10.885 3.505 11.225 4.100 ;
        RECT  9.725 0.630 12.965 0.860 ;
        RECT  12.155 0.630 12.965 0.950 ;
        RECT  9.725 0.630 10.020 1.500 ;
        RECT  10.830 1.100 11.170 1.440 ;
        RECT  10.830 1.210 12.060 1.440 ;
        RECT  11.830 1.210 12.060 3.275 ;
        RECT  12.995 2.860 14.890 3.090 ;
        RECT  14.595 2.270 14.890 3.090 ;
        RECT  8.945 3.045 13.335 3.275 ;
        RECT  8.945 3.045 9.285 3.395 ;
        RECT  11.455 3.045 11.745 3.980 ;
        RECT  12.290 1.180 14.960 1.410 ;
        RECT  14.620 1.080 14.960 1.420 ;
        RECT  12.290 1.180 12.630 1.730 ;
        RECT  14.730 1.080 14.960 2.040 ;
        RECT  14.730 1.810 15.350 2.040 ;
        RECT  15.120 2.250 17.605 2.480 ;
        RECT  17.265 2.250 17.605 2.590 ;
        RECT  15.120 1.810 15.350 3.550 ;
        RECT  14.315 3.320 15.350 3.550 ;
        RECT  14.315 3.320 14.655 3.660 ;
        RECT  1.375 1.860 3.30 2.095 ;
        RECT  0.965 1.355 3.70 1.585 ;
        RECT  2.840 3.045 3.30 3.275 ;
        RECT  2.030 3.505 3.70 3.735 ;
        RECT  0.180 3.600 1.10 3.830 ;
        RECT  4.120 0.630 5.30 0.860 ;
        RECT  1.795 0.895 3.20 1.125 ;
        RECT  7.255 2.450 10.80 2.680 ;
        RECT  9.725 0.630 11.60 0.860 ;
        RECT  8.945 3.045 12.60 3.275 ;
        RECT  12.290 1.180 13.90 1.410 ;
        RECT  15.120 2.250 16.80 2.480 ;
    END
END DFRRSX4

MACRO DFRRSX2
    CLASS CORE ;
    FOREIGN DFRRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 1.240 15.010 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.350 2.860 14.365 3.090 ;
        RECT  14.135 0.950 14.365 3.090 ;
        RECT  13.350 0.950 14.365 1.180 ;
        RECT  13.350 2.860 13.735 4.180 ;
        RECT  13.350 0.820 13.690 1.180 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.790 1.920 11.215 2.630 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.075 6.920 2.630 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.445 1.640 11.915 2.160 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.850 1.640 5.190 2.100 ;
        RECT  4.535 1.640 5.190 2.020 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  14.110 3.950 15.570 5.280 ;
        RECT  12.630 3.785 12.970 5.280 ;
        RECT  11.190 3.730 11.530 5.280 ;
        RECT  10.200 3.860 10.540 5.280 ;
        RECT  7.730 3.480 8.070 5.280 ;
        RECT  6.430 3.525 6.770 5.280 ;
        RECT  5.130 3.525 5.470 5.280 ;
        RECT  1.500 3.805 2.900 5.280 ;
        RECT  0.180 3.780 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  14.110 -0.400 15.570 0.720 ;
        RECT  12.590 -0.400 12.930 0.720 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  6.060 -0.400 6.400 0.925 ;
        RECT  1.210 -0.400 1.550 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.360 0.520 2.070 ;
        RECT  0.130 1.840 2.405 2.070 ;
        RECT  2.120 1.840 2.405 2.490 ;
        RECT  0.130 1.360 0.360 3.160 ;
        RECT  0.130 2.870 1.080 3.160 ;
        RECT  2.635 1.090 3.540 1.325 ;
        RECT  0.590 2.300 0.930 2.640 ;
        RECT  0.590 2.410 1.630 2.640 ;
        RECT  1.400 2.410 1.630 3.190 ;
        RECT  1.400 2.850 2.865 3.190 ;
        RECT  2.635 1.090 2.865 3.575 ;
        RECT  2.635 3.345 3.930 3.575 ;
        RECT  3.590 3.345 3.930 3.820 ;
        RECT  1.970 0.630 4.940 0.860 ;
        RECT  4.600 0.630 4.940 1.375 ;
        RECT  1.970 0.630 2.310 1.530 ;
        RECT  7.090 1.240 7.380 1.845 ;
        RECT  5.880 1.615 7.380 1.845 ;
        RECT  5.880 1.615 6.195 2.100 ;
        RECT  7.150 1.240 7.380 3.295 ;
        RECT  7.150 2.320 8.865 2.550 ;
        RECT  8.525 2.320 8.865 2.660 ;
        RECT  3.510 2.310 3.845 3.115 ;
        RECT  3.510 2.885 5.120 3.115 ;
        RECT  7.150 2.320 7.530 3.295 ;
        RECT  4.890 3.065 7.530 3.295 ;
        RECT  6.630 0.780 7.840 1.010 ;
        RECT  6.630 0.780 6.860 1.385 ;
        RECT  5.300 1.155 6.860 1.385 ;
        RECT  5.300 1.070 5.640 1.410 ;
        RECT  7.610 0.780 7.840 1.940 ;
        RECT  3.095 1.555 4.305 1.895 ;
        RECT  7.610 1.710 8.385 1.940 ;
        RECT  8.045 1.820 9.325 2.050 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 4.520 2.655 ;
        RECT  5.420 1.155 5.650 2.835 ;
        RECT  4.075 2.425 5.650 2.655 ;
        RECT  9.095 1.820 9.325 3.090 ;
        RECT  5.420 2.550 6.010 2.835 ;
        RECT  9.095 2.750 9.590 3.090 ;
        RECT  8.070 0.630 10.735 0.860 ;
        RECT  8.070 0.630 8.355 0.970 ;
        RECT  10.395 0.630 10.735 1.015 ;
        RECT  10.395 0.630 10.725 1.030 ;
        RECT  9.165 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  9.820 2.860 12.650 3.090 ;
        RECT  12.310 2.750 12.650 3.095 ;
        RECT  10.760 2.860 12.650 3.095 ;
        RECT  10.760 2.860 11.100 3.200 ;
        RECT  9.820 1.970 10.050 3.550 ;
        RECT  8.970 3.320 10.050 3.550 ;
        RECT  8.970 3.320 9.310 3.660 ;
        RECT  10.900 1.180 12.930 1.410 ;
        RECT  10.115 1.400 11.130 1.630 ;
        RECT  10.115 1.400 10.455 1.740 ;
        RECT  12.590 1.180 12.930 1.980 ;
        RECT  12.890 2.120 13.905 2.460 ;
        RECT  12.890 1.695 13.120 3.555 ;
        RECT  11.910 3.325 13.120 3.555 ;
        RECT  11.910 3.325 12.250 4.070 ;
        RECT  0.130 1.840 1.20 2.070 ;
        RECT  1.970 0.630 3.80 0.860 ;
        RECT  4.890 3.065 6.30 3.295 ;
        RECT  8.070 0.630 9.70 0.860 ;
        RECT  9.820 2.860 11.30 3.090 ;
        RECT  10.900 1.180 11.70 1.410 ;
    END
END DFRRSX2

MACRO DFRRSX1
    CLASS CORE ;
    FOREIGN DFRRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.285 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.640 11.845 2.305 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.835 2.045 11.215 2.630 ;
        RECT  10.520 2.045 11.215 2.385 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.585 2.075 7.120 2.360 ;
        RECT  6.425 2.250 6.805 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.710  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 2.250 13.735 2.630 ;
        RECT  12.790 2.870 13.585 3.100 ;
        RECT  13.355 1.235 13.585 3.100 ;
        RECT  12.640 1.235 13.585 1.465 ;
        RECT  12.530 3.635 13.020 3.920 ;
        RECT  12.790 2.870 13.020 3.920 ;
        RECT  12.640 0.700 12.870 1.465 ;
        RECT  12.530 0.700 12.870 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 3.270 14.365 4.180 ;
        RECT  13.970 0.820 14.310 1.160 ;
        RECT  13.970 0.820 14.200 4.180 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.250 -0.400 13.590 1.005 ;
        RECT  11.275 -0.400 11.615 0.880 ;
        RECT  6.295 -0.400 6.635 0.925 ;
        RECT  1.210 -0.400 1.550 1.450 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.250 3.330 13.590 5.280 ;
        RECT  11.990 4.170 12.330 5.280 ;
        RECT  10.415 3.665 10.755 5.280 ;
        RECT  7.815 3.480 8.155 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.215 ;
        RECT  0.170 1.985 2.445 2.215 ;
        RECT  2.160 1.985 2.445 2.325 ;
        RECT  0.170 0.645 0.400 3.360 ;
        RECT  0.170 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 0.970 2.785 ;
        RECT  0.630 2.520 1.985 2.785 ;
        RECT  1.755 2.520 1.985 3.340 ;
        RECT  1.755 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  1.970 0.630 5.135 0.860 ;
        RECT  4.795 0.630 5.135 1.280 ;
        RECT  1.970 0.630 2.310 1.450 ;
        RECT  7.325 1.240 7.665 1.845 ;
        RECT  5.975 1.615 7.665 1.845 ;
        RECT  5.975 1.615 6.255 2.095 ;
        RECT  5.975 1.615 6.235 2.120 ;
        RECT  7.380 1.240 7.665 2.690 ;
        RECT  7.380 2.460 8.830 2.690 ;
        RECT  8.490 2.460 8.830 2.800 ;
        RECT  3.520 2.285 3.845 3.115 ;
        RECT  7.265 2.720 7.615 3.295 ;
        RECT  3.520 2.885 5.120 3.115 ;
        RECT  7.380 1.240 7.615 3.295 ;
        RECT  4.890 3.065 7.615 3.295 ;
        RECT  6.865 0.780 8.125 1.010 ;
        RECT  5.515 1.070 5.875 1.385 ;
        RECT  6.865 0.780 7.095 1.385 ;
        RECT  5.515 1.155 7.095 1.385 ;
        RECT  5.515 1.070 5.870 1.410 ;
        RECT  3.135 1.555 4.305 1.785 ;
        RECT  7.895 0.780 8.125 2.020 ;
        RECT  3.135 1.555 3.420 1.895 ;
        RECT  7.895 1.790 9.290 2.020 ;
        RECT  8.775 1.790 9.290 2.130 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 4.550 2.655 ;
        RECT  4.075 2.425 5.745 2.655 ;
        RECT  5.515 1.070 5.745 2.655 ;
        RECT  5.535 2.550 6.040 2.835 ;
        RECT  9.060 1.790 9.290 3.240 ;
        RECT  9.060 2.900 9.590 3.240 ;
        RECT  8.355 0.630 10.810 0.860 ;
        RECT  10.470 0.630 10.810 0.950 ;
        RECT  8.355 0.630 8.695 0.970 ;
        RECT  9.135 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  9.625 1.970 10.150 2.200 ;
        RECT  11.470 2.635 12.050 2.945 ;
        RECT  9.920 2.860 11.700 3.200 ;
        RECT  9.920 1.970 10.150 3.710 ;
        RECT  8.970 3.480 10.150 3.710 ;
        RECT  8.970 3.480 9.310 3.820 ;
        RECT  10.085 1.180 12.340 1.410 ;
        RECT  10.085 1.180 10.425 1.720 ;
        RECT  12.110 1.180 12.340 1.925 ;
        RECT  12.330 1.695 12.900 2.500 ;
        RECT  12.330 2.160 13.050 2.500 ;
        RECT  12.330 1.695 12.560 3.405 ;
        RECT  12.030 3.175 12.560 3.405 ;
        RECT  12.030 3.175 12.260 3.895 ;
        RECT  11.190 3.665 12.260 3.895 ;
        RECT  11.190 3.665 11.530 4.005 ;
        RECT  0.170 1.985 1.90 2.215 ;
        RECT  1.970 0.630 4.70 0.860 ;
        RECT  4.890 3.065 6.80 3.295 ;
        RECT  8.355 0.630 9.30 0.860 ;
        RECT  10.085 1.180 11.20 1.410 ;
    END
END DFRRSX1

MACRO DFRRSX0
    CLASS CORE ;
    FOREIGN DFRRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.260 2.135 6.805 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.592  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.065 2.860 12.625 3.350 ;
        RECT  12.395 0.630 12.625 3.350 ;
        RECT  11.730 0.630 12.625 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.380 2.235 4.915 2.695 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.250 10.220 2.760 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.248  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.660 2.250 11.215 2.845 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.443  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.855 3.010 13.735 3.350 ;
        RECT  13.335 2.860 13.735 3.350 ;
        RECT  13.335 1.170 13.565 3.350 ;
        RECT  12.855 1.170 13.565 1.510 ;
        END
    END QN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.120 3.810 13.040 5.280 ;
        RECT  9.565 3.910 9.900 5.280 ;
        RECT  6.970 3.630 7.310 5.280 ;
        RECT  4.810 3.910 6.085 5.280 ;
        RECT  1.470 3.520 2.335 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.865 -0.400 13.205 0.710 ;
        RECT  10.700 -0.400 11.040 0.950 ;
        RECT  6.030 -0.400 6.315 1.400 ;
        RECT  1.100 -0.400 1.440 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.970 ;
        RECT  0.115 1.740 2.335 1.970 ;
        RECT  2.050 1.740 2.335 2.460 ;
        RECT  0.115 0.630 0.345 3.060 ;
        RECT  0.115 2.770 1.010 3.060 ;
        RECT  2.565 1.285 3.470 1.545 ;
        RECT  0.575 2.200 1.565 2.540 ;
        RECT  1.335 2.200 1.565 3.060 ;
        RECT  1.335 2.690 2.795 3.060 ;
        RECT  2.565 1.285 2.795 4.140 ;
        RECT  2.565 3.910 3.810 4.140 ;
        RECT  3.470 3.910 3.810 4.250 ;
        RECT  1.900 0.825 4.870 1.055 ;
        RECT  1.900 0.825 2.240 1.510 ;
        RECT  4.530 0.825 4.870 1.545 ;
        RECT  7.005 1.230 7.265 1.570 ;
        RECT  5.605 2.160 5.945 2.500 ;
        RECT  7.035 1.230 7.265 3.200 ;
        RECT  3.190 2.840 3.530 3.180 ;
        RECT  5.715 2.860 8.260 3.200 ;
        RECT  3.300 2.840 3.530 3.675 ;
        RECT  5.715 2.160 5.945 3.675 ;
        RECT  3.300 3.445 5.945 3.675 ;
        RECT  6.545 0.765 7.725 0.995 ;
        RECT  5.145 1.230 5.570 1.905 ;
        RECT  5.145 1.675 6.775 1.905 ;
        RECT  6.545 0.765 6.775 1.905 ;
        RECT  3.025 1.775 5.375 2.005 ;
        RECT  3.025 1.775 4.090 2.180 ;
        RECT  7.495 0.765 7.725 2.485 ;
        RECT  7.495 2.190 8.875 2.485 ;
        RECT  3.860 1.775 4.090 3.180 ;
        RECT  5.145 1.230 5.375 3.200 ;
        RECT  3.860 2.840 4.200 3.180 ;
        RECT  5.145 2.860 5.485 3.200 ;
        RECT  8.590 2.190 8.875 3.435 ;
        RECT  7.955 0.630 10.170 0.860 ;
        RECT  7.955 0.630 8.240 0.970 ;
        RECT  9.830 0.630 10.170 0.970 ;
        RECT  8.800 1.170 9.140 1.510 ;
        RECT  10.140 3.075 10.500 3.525 ;
        RECT  10.140 3.125 11.375 3.525 ;
        RECT  9.105 3.285 11.375 3.525 ;
        RECT  9.105 1.280 9.335 3.970 ;
        RECT  8.270 3.665 9.335 3.970 ;
        RECT  11.730 1.310 12.070 2.170 ;
        RECT  9.750 1.690 12.070 1.920 ;
        RECT  9.750 1.690 10.090 2.020 ;
        RECT  11.605 1.830 12.165 2.170 ;
        RECT  11.605 1.690 11.835 4.155 ;
        RECT  10.695 3.925 11.835 4.155 ;
        RECT  10.695 3.925 11.035 4.250 ;
        RECT  0.115 1.740 1.80 1.970 ;
        RECT  1.900 0.825 3.60 1.055 ;
        RECT  5.715 2.860 7.40 3.200 ;
        RECT  3.300 3.445 4.90 3.675 ;
        RECT  3.025 1.775 4.40 2.005 ;
        RECT  7.955 0.630 9.60 0.860 ;
        RECT  9.105 3.285 10.50 3.525 ;
        RECT  9.750 1.690 11.30 1.920 ;
    END
END DFRRSX0

MACRO DFRRSQX4
    CLASS CORE ;
    FOREIGN DFRRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 1.240 17.460 4.030 ;
        RECT  15.800 2.250 17.460 2.630 ;
        RECT  15.800 0.790 16.140 2.630 ;
        RECT  15.680 2.790 16.030 4.030 ;
        RECT  15.800 0.790 16.030 4.030 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.905 1.640 14.365 2.560 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.655 2.230 13.265 2.630 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.685 1.660 8.495 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.560 -0.400 16.900 0.720 ;
        RECT  15.040 -0.400 15.380 0.835 ;
        RECT  13.430 -0.400 13.770 0.710 ;
        RECT  7.830 -0.400 8.115 0.970 ;
        RECT  2.255 -0.400 3.825 0.665 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.400 2.860 16.740 5.280 ;
        RECT  14.875 4.060 15.215 5.280 ;
        RECT  12.435 3.910 13.895 5.280 ;
        RECT  10.135 3.965 10.475 5.280 ;
        RECT  7.715 2.910 8.015 5.280 ;
        RECT  2.410 3.965 3.845 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.765 1.815 2.105 2.095 ;
        RECT  1.375 1.860 4.020 2.095 ;
        RECT  3.790 1.860 4.020 2.800 ;
        RECT  3.790 2.460 4.130 2.800 ;
        RECT  1.375 1.860 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.965 1.355 4.535 1.585 ;
        RECT  0.965 1.290 1.305 1.630 ;
        RECT  2.925 1.355 4.535 1.630 ;
        RECT  4.245 1.355 4.535 1.695 ;
        RECT  5.475 1.160 5.810 1.500 ;
        RECT  4.765 1.270 5.810 1.500 ;
        RECT  1.835 2.325 3.180 2.665 ;
        RECT  2.840 2.325 3.180 3.275 ;
        RECT  4.765 1.270 4.995 3.540 ;
        RECT  2.840 3.045 4.995 3.275 ;
        RECT  4.735 3.200 5.080 3.540 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.415 3.735 ;
        RECT  4.185 3.505 4.415 4.000 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  5.500 2.980 5.840 4.000 ;
        RECT  4.185 3.770 5.840 4.000 ;
        RECT  0.365 0.640 0.705 1.015 ;
        RECT  4.120 0.630 6.270 0.860 ;
        RECT  1.375 1.860 3.40 2.095 ;
        RECT  0.965 1.355 3.60 1.585 ;
        RECT  2.840 3.045 3.50 3.275 ;
        RECT  2.030 3.505 3.20 3.735 ;
        RECT  0.180 3.600 1.60 3.830 ;
        RECT  4.120 0.630 5.40 0.860 ;
        RECT  0.365 0.785 2.025 1.015 ;
        RECT  4.120 0.630 4.350 1.125 ;
        RECT  1.795 0.895 4.350 1.125 ;
        RECT  6.040 0.630 6.270 1.660 ;
        RECT  6.040 1.320 6.625 1.660 ;
        RECT  8.345 0.775 9.495 1.005 ;
        RECT  6.500 0.735 7.370 1.090 ;
        RECT  8.345 0.775 8.575 1.430 ;
        RECT  7.140 1.200 8.575 1.430 ;
        RECT  9.265 0.775 9.495 2.090 ;
        RECT  9.265 1.860 10.930 2.090 ;
        RECT  7.140 0.735 7.370 2.150 ;
        RECT  6.740 1.920 7.370 2.150 ;
        RECT  10.590 1.860 10.930 2.200 ;
        RECT  6.740 1.920 7.025 3.195 ;
        RECT  5.225 1.820 5.535 2.175 ;
        RECT  11.260 1.670 11.600 2.010 ;
        RECT  5.225 1.945 6.510 2.175 ;
        RECT  8.805 1.240 9.035 2.680 ;
        RECT  8.805 2.340 9.505 2.680 ;
        RECT  11.260 1.670 11.490 2.680 ;
        RECT  7.255 2.450 11.490 2.680 ;
        RECT  8.395 2.450 8.735 2.860 ;
        RECT  6.170 1.945 6.510 3.655 ;
        RECT  8.395 2.450 8.625 3.855 ;
        RECT  7.255 2.450 7.485 3.655 ;
        RECT  6.170 3.425 7.485 3.655 ;
        RECT  9.605 3.505 11.115 3.735 ;
        RECT  10.885 3.505 11.115 4.100 ;
        RECT  8.395 3.625 9.835 3.855 ;
        RECT  10.885 3.760 11.225 4.100 ;
        RECT  9.725 0.630 12.965 0.860 ;
        RECT  12.155 0.630 12.965 0.950 ;
        RECT  9.725 0.630 10.020 1.500 ;
        RECT  10.830 1.100 11.170 1.440 ;
        RECT  10.830 1.210 12.060 1.440 ;
        RECT  11.830 1.210 12.060 3.275 ;
        RECT  12.995 2.860 14.890 3.090 ;
        RECT  14.595 2.270 14.890 3.090 ;
        RECT  8.945 3.045 13.335 3.275 ;
        RECT  8.945 3.045 9.285 3.395 ;
        RECT  11.455 3.045 11.745 3.980 ;
        RECT  14.415 1.110 14.825 1.410 ;
        RECT  12.290 1.180 14.825 1.410 ;
        RECT  14.435 1.110 14.825 1.420 ;
        RECT  12.290 1.180 12.630 1.675 ;
        RECT  14.595 1.110 14.825 2.040 ;
        RECT  14.595 1.810 15.350 2.040 ;
        RECT  15.120 1.810 15.350 3.550 ;
        RECT  14.315 3.320 15.350 3.550 ;
        RECT  14.315 3.320 14.655 3.660 ;
    END
END DFRRSQX4

MACRO DFRRSQX2
    CLASS CORE ;
    FOREIGN DFRRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 1.240 13.750 3.550 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.780 2.070 11.225 2.630 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.075 6.920 2.630 ;
        END
    END C
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.640 11.845 2.585 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.850 1.640 5.190 2.100 ;
        RECT  4.535 1.640 5.190 2.020 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  12.850 3.950 14.310 5.280 ;
        RECT  11.370 3.730 11.710 5.280 ;
        RECT  10.000 3.910 10.340 5.280 ;
        RECT  7.730 3.480 8.070 5.280 ;
        RECT  6.430 3.525 6.770 5.280 ;
        RECT  5.130 3.525 5.470 5.280 ;
        RECT  1.500 3.805 2.900 5.280 ;
        RECT  0.180 3.780 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  12.850 -0.400 14.310 0.720 ;
        RECT  11.155 -0.400 11.495 0.950 ;
        RECT  6.060 -0.400 6.400 0.925 ;
        RECT  1.210 -0.400 1.550 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.360 0.520 2.070 ;
        RECT  0.130 1.840 2.405 2.070 ;
        RECT  2.120 1.840 2.405 2.490 ;
        RECT  0.130 1.360 0.360 3.100 ;
        RECT  0.130 2.870 1.080 3.100 ;
        RECT  0.740 2.870 1.080 3.160 ;
        RECT  2.635 1.090 3.540 1.325 ;
        RECT  0.590 2.300 0.930 2.640 ;
        RECT  0.590 2.410 1.630 2.640 ;
        RECT  1.400 2.410 1.630 3.190 ;
        RECT  1.400 2.850 2.865 3.190 ;
        RECT  2.635 1.090 2.865 3.575 ;
        RECT  2.635 3.345 3.930 3.575 ;
        RECT  3.590 3.345 3.930 3.820 ;
        RECT  1.970 0.630 4.940 0.860 ;
        RECT  4.600 0.630 4.940 1.375 ;
        RECT  1.970 0.630 2.310 1.530 ;
        RECT  7.090 1.240 7.380 1.845 ;
        RECT  5.880 1.615 7.380 1.845 ;
        RECT  5.880 1.615 6.195 2.100 ;
        RECT  7.150 1.240 7.380 3.295 ;
        RECT  7.150 2.320 8.865 2.550 ;
        RECT  8.525 2.320 8.865 2.660 ;
        RECT  3.510 2.310 3.845 3.115 ;
        RECT  3.510 2.885 5.120 3.115 ;
        RECT  7.150 2.320 7.530 3.295 ;
        RECT  4.890 3.065 7.530 3.295 ;
        RECT  6.630 0.780 7.840 1.010 ;
        RECT  6.630 0.780 6.860 1.385 ;
        RECT  5.300 1.155 6.860 1.385 ;
        RECT  5.300 1.070 5.640 1.410 ;
        RECT  3.095 1.555 3.390 1.895 ;
        RECT  7.610 0.780 7.840 1.940 ;
        RECT  3.095 1.665 4.305 1.895 ;
        RECT  7.610 1.710 8.385 1.940 ;
        RECT  8.045 1.820 9.325 2.050 ;
        RECT  4.075 1.665 4.305 2.655 ;
        RECT  4.075 2.290 4.520 2.655 ;
        RECT  5.420 1.155 5.650 2.835 ;
        RECT  4.075 2.425 5.650 2.655 ;
        RECT  9.095 1.820 9.325 3.080 ;
        RECT  5.420 2.550 6.010 2.835 ;
        RECT  9.095 2.740 9.590 3.080 ;
        RECT  8.070 0.630 10.735 0.860 ;
        RECT  8.070 0.630 8.355 0.970 ;
        RECT  10.395 0.630 10.735 1.040 ;
        RECT  9.165 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  12.320 2.750 12.660 3.090 ;
        RECT  9.820 2.860 12.660 3.090 ;
        RECT  10.760 2.860 11.100 3.200 ;
        RECT  9.820 1.970 10.050 3.550 ;
        RECT  8.950 3.320 10.050 3.550 ;
        RECT  8.950 3.320 9.290 3.660 ;
        RECT  11.985 0.630 12.325 1.410 ;
        RECT  10.985 1.180 13.120 1.410 ;
        RECT  10.115 1.400 11.215 1.630 ;
        RECT  10.115 1.400 10.455 1.740 ;
        RECT  12.890 1.180 13.120 3.720 ;
        RECT  12.090 3.490 13.120 3.720 ;
        RECT  12.090 3.490 12.430 4.060 ;
        RECT  0.130 1.840 1.80 2.070 ;
        RECT  1.970 0.630 3.80 0.860 ;
        RECT  4.890 3.065 6.70 3.295 ;
        RECT  8.070 0.630 9.00 0.860 ;
        RECT  9.820 2.860 11.60 3.090 ;
        RECT  10.985 1.180 12.50 1.410 ;
    END
END DFRRSQX2

MACRO DFRRSQX1
    CLASS CORE ;
    FOREIGN DFRRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.285 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.640 11.845 2.305 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.835 2.045 11.215 2.630 ;
        RECT  10.520 2.045 11.215 2.385 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.585 2.075 7.120 2.360 ;
        RECT  6.425 2.250 6.805 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.712  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.880 2.400 13.735 2.630 ;
        RECT  13.355 2.250 13.735 2.630 ;
        RECT  13.355 1.235 13.585 2.630 ;
        RECT  12.730 1.235 13.585 1.465 ;
        RECT  12.620 3.635 13.110 3.920 ;
        RECT  12.880 2.400 13.110 3.920 ;
        RECT  12.730 0.700 12.960 1.465 ;
        RECT  12.655 3.615 13.110 3.920 ;
        RECT  12.620 0.700 12.960 1.040 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.340 -0.400 13.680 1.005 ;
        RECT  11.275 -0.400 11.615 0.870 ;
        RECT  6.295 -0.400 6.635 0.925 ;
        RECT  1.210 -0.400 1.550 1.450 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  13.340 3.330 13.680 5.280 ;
        RECT  11.990 4.170 12.330 5.280 ;
        RECT  10.415 3.665 10.755 5.280 ;
        RECT  7.815 3.480 8.155 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.215 ;
        RECT  0.170 1.985 2.445 2.215 ;
        RECT  2.160 1.985 2.445 2.325 ;
        RECT  0.170 0.645 0.400 3.360 ;
        RECT  0.170 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 0.970 2.785 ;
        RECT  0.630 2.520 1.985 2.785 ;
        RECT  1.755 2.520 1.985 3.340 ;
        RECT  1.755 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  1.970 0.630 5.135 0.860 ;
        RECT  4.795 0.630 5.135 1.280 ;
        RECT  1.970 0.630 2.310 1.450 ;
        RECT  7.325 1.240 7.665 1.845 ;
        RECT  5.975 1.615 7.665 1.845 ;
        RECT  5.975 1.615 6.255 2.095 ;
        RECT  5.975 1.615 6.235 2.120 ;
        RECT  7.380 1.240 7.665 2.690 ;
        RECT  7.380 2.460 8.830 2.690 ;
        RECT  8.490 2.460 8.830 2.800 ;
        RECT  3.520 2.305 3.845 3.115 ;
        RECT  7.265 2.720 7.615 3.295 ;
        RECT  3.520 2.885 5.120 3.115 ;
        RECT  7.380 1.240 7.615 3.295 ;
        RECT  4.890 3.065 7.615 3.295 ;
        RECT  6.865 0.780 8.125 1.010 ;
        RECT  5.515 1.070 5.875 1.385 ;
        RECT  6.865 0.780 7.095 1.385 ;
        RECT  5.515 1.155 7.095 1.385 ;
        RECT  5.515 1.070 5.870 1.410 ;
        RECT  3.135 1.555 4.305 1.785 ;
        RECT  7.895 0.780 8.125 2.020 ;
        RECT  3.135 1.555 3.420 1.895 ;
        RECT  7.895 1.790 9.290 2.020 ;
        RECT  8.805 1.790 9.290 2.130 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 4.550 2.655 ;
        RECT  4.075 2.425 5.745 2.655 ;
        RECT  5.515 1.070 5.745 2.655 ;
        RECT  5.535 2.550 6.040 2.835 ;
        RECT  9.060 1.790 9.290 3.130 ;
        RECT  9.250 2.900 9.590 3.240 ;
        RECT  8.355 0.630 10.810 0.860 ;
        RECT  10.470 0.630 10.810 0.950 ;
        RECT  8.355 0.630 8.695 0.970 ;
        RECT  9.135 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  9.625 1.970 10.150 2.200 ;
        RECT  11.470 2.635 12.050 2.945 ;
        RECT  9.920 2.860 11.700 3.200 ;
        RECT  9.920 1.970 10.150 3.710 ;
        RECT  8.970 3.480 10.150 3.710 ;
        RECT  8.970 3.480 9.310 3.820 ;
        RECT  10.085 1.180 12.340 1.410 ;
        RECT  10.085 1.180 10.425 1.730 ;
        RECT  12.110 1.180 12.340 1.925 ;
        RECT  12.330 1.695 12.910 1.980 ;
        RECT  12.330 1.695 12.560 3.405 ;
        RECT  12.030 3.175 12.560 3.405 ;
        RECT  12.030 3.175 12.260 3.895 ;
        RECT  11.190 3.665 12.260 3.895 ;
        RECT  11.190 3.665 11.530 4.005 ;
        RECT  0.170 1.985 1.60 2.215 ;
        RECT  1.970 0.630 4.60 0.860 ;
        RECT  4.890 3.065 6.30 3.295 ;
        RECT  8.355 0.630 9.20 0.860 ;
        RECT  10.085 1.180 11.40 1.410 ;
    END
END DFRRSQX1

MACRO DFRRSQX0
    CLASS CORE ;
    FOREIGN DFRRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.260 2.135 6.805 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.592  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.065 2.860 12.485 3.350 ;
        RECT  12.255 0.630 12.485 3.350 ;
        RECT  11.730 0.630 12.485 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.380 2.235 4.915 2.695 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.250 10.220 2.760 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.248  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.660 2.250 11.215 2.845 ;
        END
    END SN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  12.065 3.810 12.405 5.280 ;
        RECT  9.565 3.910 9.900 5.280 ;
        RECT  6.970 3.630 7.310 5.280 ;
        RECT  4.810 3.910 6.085 5.280 ;
        RECT  1.470 3.520 2.335 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.700 -0.400 11.040 0.950 ;
        RECT  6.030 -0.400 6.315 1.400 ;
        RECT  1.100 -0.400 1.440 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.970 ;
        RECT  0.115 1.740 2.335 1.970 ;
        RECT  2.050 1.740 2.335 2.460 ;
        RECT  0.115 0.630 0.345 3.060 ;
        RECT  0.115 2.770 1.010 3.060 ;
        RECT  2.565 1.285 3.470 1.545 ;
        RECT  0.575 2.200 1.565 2.540 ;
        RECT  1.335 2.200 1.565 3.060 ;
        RECT  1.335 2.690 2.795 3.060 ;
        RECT  2.565 1.285 2.795 4.140 ;
        RECT  2.565 3.910 3.810 4.140 ;
        RECT  3.470 3.910 3.810 4.250 ;
        RECT  1.900 0.825 4.870 1.055 ;
        RECT  1.900 0.825 2.240 1.510 ;
        RECT  4.530 0.825 4.870 1.545 ;
        RECT  7.005 1.230 7.265 1.570 ;
        RECT  5.605 2.160 5.945 2.500 ;
        RECT  7.035 1.230 7.265 3.200 ;
        RECT  3.190 2.840 3.530 3.180 ;
        RECT  5.715 2.860 8.260 3.200 ;
        RECT  3.300 2.840 3.530 3.675 ;
        RECT  5.715 2.160 5.945 3.675 ;
        RECT  3.300 3.445 5.945 3.675 ;
        RECT  6.545 0.765 7.725 0.995 ;
        RECT  5.145 1.230 5.570 1.905 ;
        RECT  5.145 1.675 6.775 1.905 ;
        RECT  6.545 0.765 6.775 1.905 ;
        RECT  3.025 1.775 5.375 2.005 ;
        RECT  3.025 1.775 4.090 2.180 ;
        RECT  7.495 0.765 7.725 2.485 ;
        RECT  7.495 2.190 8.875 2.485 ;
        RECT  3.860 1.775 4.090 3.180 ;
        RECT  5.145 1.230 5.375 3.200 ;
        RECT  3.860 2.840 4.200 3.180 ;
        RECT  5.145 2.860 5.485 3.200 ;
        RECT  8.590 2.190 8.875 3.435 ;
        RECT  7.955 0.630 10.170 0.860 ;
        RECT  7.955 0.630 8.240 0.970 ;
        RECT  9.830 0.630 10.170 0.970 ;
        RECT  8.800 1.170 9.140 1.510 ;
        RECT  10.140 3.075 10.500 3.525 ;
        RECT  9.105 3.125 11.375 3.525 ;
        RECT  9.105 1.280 9.335 3.970 ;
        RECT  8.270 3.665 9.335 3.970 ;
        RECT  9.750 1.310 12.025 1.540 ;
        RECT  11.605 1.310 12.025 1.650 ;
        RECT  9.750 1.310 10.090 2.020 ;
        RECT  11.605 1.310 11.835 4.155 ;
        RECT  10.695 3.925 11.835 4.155 ;
        RECT  10.695 3.925 11.035 4.250 ;
        RECT  0.115 1.740 1.80 1.970 ;
        RECT  1.900 0.825 3.40 1.055 ;
        RECT  5.715 2.860 7.90 3.200 ;
        RECT  3.300 3.445 4.50 3.675 ;
        RECT  3.025 1.775 4.60 2.005 ;
        RECT  7.955 0.630 9.80 0.860 ;
        RECT  9.105 3.125 10.50 3.525 ;
        RECT  9.750 1.310 11.70 1.540 ;
    END
END DFRRSQX0

MACRO DFRRQX4
    CLASS CORE ;
    FOREIGN DFRRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 2.075 16.885 3.880 ;
        RECT  14.330 2.075 16.885 2.305 ;
        RECT  15.770 1.130 16.110 2.305 ;
        RECT  15.050 2.075 15.390 3.880 ;
        RECT  14.330 1.130 14.670 2.305 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.290 1.640 13.105 2.020 ;
        RECT  12.290 1.640 12.630 2.190 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.055 1.660 7.850 2.225 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.760 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 1.470 ;
        RECT  15.050 -0.400 15.390 1.470 ;
        RECT  12.800 -0.400 13.140 0.950 ;
        RECT  7.230 -0.400 7.515 0.970 ;
        RECT  1.750 -0.400 3.225 0.655 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 2.640 16.110 5.280 ;
        RECT  14.330 2.640 14.670 5.280 ;
        RECT  11.490 3.760 12.950 5.280 ;
        RECT  9.315 4.170 9.655 5.280 ;
        RECT  6.825 3.925 7.165 5.280 ;
        RECT  2.410 3.985 3.245 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.805 1.920 2.090 ;
        RECT  1.375 1.860 3.420 2.090 ;
        RECT  3.190 1.860 3.420 2.800 ;
        RECT  3.190 2.460 3.530 2.800 ;
        RECT  1.375 1.805 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.780 1.345 3.935 1.575 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  2.325 1.345 3.935 1.630 ;
        RECT  3.645 1.345 3.935 1.695 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.525 5.200 3.755 ;
        RECT  4.860 3.010 5.200 3.755 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  4.875 1.160 5.210 1.500 ;
        RECT  4.165 1.270 5.210 1.500 ;
        RECT  1.835 2.325 2.580 2.665 ;
        RECT  4.165 1.270 4.395 3.295 ;
        RECT  2.240 2.325 2.580 3.295 ;
        RECT  4.140 2.955 4.480 3.295 ;
        RECT  2.240 3.065 4.480 3.295 ;
        RECT  0.180 0.640 0.520 1.015 ;
        RECT  3.520 0.700 5.670 0.930 ;
        RECT  0.180 0.785 1.520 1.015 ;
        RECT  1.290 0.885 3.750 1.115 ;
        RECT  5.440 0.700 5.670 1.655 ;
        RECT  5.440 1.315 6.025 1.655 ;
        RECT  7.745 0.775 8.895 1.005 ;
        RECT  5.900 0.735 6.770 1.085 ;
        RECT  6.255 0.735 6.770 1.430 ;
        RECT  7.745 0.775 7.975 1.430 ;
        RECT  6.255 1.200 7.975 1.430 ;
        RECT  8.665 0.775 8.895 2.090 ;
        RECT  8.665 1.860 10.330 2.090 ;
        RECT  6.255 0.735 6.485 2.150 ;
        RECT  9.990 1.860 10.330 2.200 ;
        RECT  6.050 1.920 6.390 3.235 ;
        RECT  4.625 1.820 4.935 2.175 ;
        RECT  10.660 1.670 11.000 1.980 ;
        RECT  4.625 1.945 5.810 2.175 ;
        RECT  8.205 1.240 8.435 2.805 ;
        RECT  8.205 2.340 8.685 2.805 ;
        RECT  8.205 2.520 10.890 2.805 ;
        RECT  10.660 1.670 10.890 2.805 ;
        RECT  7.585 2.575 10.890 2.805 ;
        RECT  7.585 2.575 7.925 2.915 ;
        RECT  5.470 1.945 5.810 3.695 ;
        RECT  5.470 3.465 7.815 3.695 ;
        RECT  7.585 2.575 7.815 3.940 ;
        RECT  7.585 3.710 10.170 3.940 ;
        RECT  9.940 3.710 10.170 4.250 ;
        RECT  9.940 3.965 10.280 4.250 ;
        RECT  9.125 0.630 12.340 0.860 ;
        RECT  11.530 0.630 12.340 0.950 ;
        RECT  9.125 0.630 9.420 1.500 ;
        RECT  10.230 1.100 10.570 1.440 ;
        RECT  10.230 1.210 11.460 1.440 ;
        RECT  13.295 2.150 13.600 2.650 ;
        RECT  13.315 2.120 13.600 2.650 ;
        RECT  11.230 2.420 13.600 2.650 ;
        RECT  12.050 2.420 12.390 3.150 ;
        RECT  11.230 1.210 11.460 3.395 ;
        RECT  8.125 3.165 11.460 3.395 ;
        RECT  8.125 3.165 8.465 3.480 ;
        RECT  10.485 3.165 10.800 3.860 ;
        RECT  10.510 3.165 10.800 3.890 ;
        RECT  11.690 1.180 14.060 1.410 ;
        RECT  13.560 1.180 14.060 1.520 ;
        RECT  11.690 1.180 11.975 1.730 ;
        RECT  13.830 1.180 14.060 3.240 ;
        RECT  13.570 3.010 13.910 3.880 ;
        RECT  1.375 1.860 2.70 2.090 ;
        RECT  0.780 1.345 2.30 1.575 ;
        RECT  2.030 3.525 4.20 3.755 ;
        RECT  0.180 3.600 1.60 3.830 ;
        RECT  2.240 3.065 3.80 3.295 ;
        RECT  3.520 0.700 4.90 0.930 ;
        RECT  1.290 0.885 2.50 1.115 ;
        RECT  8.205 2.520 9.60 2.805 ;
        RECT  7.585 2.575 9.70 2.805 ;
        RECT  5.470 3.465 6.60 3.695 ;
        RECT  7.585 3.710 9.90 3.940 ;
        RECT  9.125 0.630 11.70 0.860 ;
        RECT  11.230 2.420 12.60 2.650 ;
        RECT  8.125 3.165 10.70 3.395 ;
        RECT  11.690 1.180 13.60 1.410 ;
    END
END DFRRQX4

MACRO DFRRQX2
    CLASS CORE ;
    FOREIGN DFRRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 1.240 12.490 3.550 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.045 2.220 10.605 2.680 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.075 6.390 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.400 1.640 4.915 2.120 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  11.590 3.950 13.050 5.280 ;
        RECT  9.620 4.170 9.960 5.280 ;
        RECT  7.200 3.660 7.540 5.280 ;
        RECT  5.900 3.525 6.240 5.280 ;
        RECT  4.600 3.525 4.940 5.280 ;
        RECT  1.470 3.805 2.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.590 -0.400 13.050 0.720 ;
        RECT  10.230 -0.400 10.570 1.040 ;
        RECT  5.390 -0.400 5.730 0.925 ;
        RECT  0.780 -0.400 1.120 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.360 0.520 2.510 ;
        RECT  0.115 2.280 1.905 2.510 ;
        RECT  1.620 2.280 1.905 2.620 ;
        RECT  0.115 2.280 0.345 4.070 ;
        RECT  0.115 3.730 0.620 4.070 ;
        RECT  2.135 1.305 3.040 1.645 ;
        RECT  0.575 2.850 2.365 3.190 ;
        RECT  2.135 1.305 2.365 3.575 ;
        RECT  2.135 3.345 3.630 3.575 ;
        RECT  3.290 3.345 3.630 3.685 ;
        RECT  1.580 0.630 4.240 0.950 ;
        RECT  1.580 0.630 1.920 1.090 ;
        RECT  6.420 1.240 6.710 1.845 ;
        RECT  5.145 1.615 6.850 1.845 ;
        RECT  5.145 1.615 5.450 2.195 ;
        RECT  6.620 1.615 6.850 3.295 ;
        RECT  7.920 2.360 8.260 2.700 ;
        RECT  6.620 2.470 8.260 2.700 ;
        RECT  3.010 2.505 3.350 3.115 ;
        RECT  3.010 2.885 4.910 3.115 ;
        RECT  6.620 2.470 7.000 3.295 ;
        RECT  4.680 3.065 7.000 3.295 ;
        RECT  5.960 0.780 7.310 1.010 ;
        RECT  4.630 1.155 6.190 1.385 ;
        RECT  5.960 0.780 6.190 1.385 ;
        RECT  4.630 1.070 4.970 1.410 ;
        RECT  3.680 1.180 4.970 1.410 ;
        RECT  7.080 0.780 7.310 1.980 ;
        RECT  7.080 1.750 7.660 1.980 ;
        RECT  7.320 1.900 8.740 2.130 ;
        RECT  2.595 1.880 3.910 2.220 ;
        RECT  3.680 1.180 3.910 2.655 ;
        RECT  3.680 2.315 4.020 2.655 ;
        RECT  3.680 2.425 5.480 2.655 ;
        RECT  8.510 1.900 8.740 3.130 ;
        RECT  5.140 2.425 5.480 2.835 ;
        RECT  8.510 2.805 9.010 3.130 ;
        RECT  7.540 0.630 9.810 0.970 ;
        RECT  9.470 0.630 9.810 1.040 ;
        RECT  8.440 1.330 9.200 1.670 ;
        RECT  8.970 1.330 9.200 2.575 ;
        RECT  8.970 2.345 9.470 2.575 ;
        RECT  9.240 2.915 11.135 3.145 ;
        RECT  10.180 2.915 11.135 3.260 ;
        RECT  10.180 2.915 10.520 3.440 ;
        RECT  9.240 2.345 9.470 3.715 ;
        RECT  8.385 3.485 9.470 3.715 ;
        RECT  8.385 3.485 8.725 3.825 ;
        RECT  10.795 1.360 11.135 1.990 ;
        RECT  9.430 1.760 11.595 1.990 ;
        RECT  9.430 1.760 9.770 2.115 ;
        RECT  11.365 1.760 11.595 3.720 ;
        RECT  10.940 3.490 11.595 3.720 ;
        RECT  10.940 3.490 11.170 4.180 ;
        RECT  10.830 3.840 11.170 4.180 ;
        RECT  1.580 0.630 3.80 0.950 ;
        RECT  4.680 3.065 6.30 3.295 ;
        RECT  7.540 0.630 8.40 0.970 ;
        RECT  9.430 1.760 10.60 1.990 ;
    END
END DFRRQX2

MACRO DFRRQX1
    CLASS CORE ;
    FOREIGN DFRRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.655 2.025 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.955 2.075 6.490 2.360 ;
        RECT  5.795 2.250 6.175 2.630 ;
        END
    END C
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.050 1.640 10.610 2.085 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.680  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.620 2.400 12.475 2.630 ;
        RECT  11.905 2.250 12.475 2.630 ;
        RECT  11.905 1.235 12.135 2.630 ;
        RECT  11.360 1.235 12.135 1.465 ;
        RECT  11.360 3.435 11.850 3.720 ;
        RECT  11.620 2.400 11.850 3.720 ;
        RECT  11.360 0.700 11.700 1.465 ;
        RECT  11.395 3.415 11.850 3.720 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.080 -0.400 12.420 1.005 ;
        RECT  10.540 -0.400 10.880 0.950 ;
        RECT  5.725 -0.400 6.065 0.925 ;
        RECT  0.915 -0.400 1.255 1.395 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  12.080 3.330 12.420 5.280 ;
        RECT  9.800 3.840 10.140 5.280 ;
        RECT  7.185 3.480 7.525 5.280 ;
        RECT  5.885 3.525 6.225 5.280 ;
        RECT  4.585 3.525 4.925 5.280 ;
        RECT  1.940 3.840 2.280 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.645 0.555 0.985 ;
        RECT  0.115 0.645 0.400 2.350 ;
        RECT  0.115 2.120 1.950 2.350 ;
        RECT  1.665 2.120 1.950 2.460 ;
        RECT  0.115 0.645 0.345 3.790 ;
        RECT  0.115 3.450 0.760 3.790 ;
        RECT  2.180 1.090 3.205 1.325 ;
        RECT  0.575 2.855 0.905 3.195 ;
        RECT  0.575 2.930 1.450 3.195 ;
        RECT  1.220 2.930 1.450 4.180 ;
        RECT  2.180 1.090 2.410 3.575 ;
        RECT  1.220 3.345 3.525 3.575 ;
        RECT  3.185 3.345 3.525 3.665 ;
        RECT  1.220 3.345 1.560 4.180 ;
        RECT  1.635 0.630 4.605 0.860 ;
        RECT  4.265 0.630 4.605 1.375 ;
        RECT  1.635 0.630 1.950 1.450 ;
        RECT  5.345 1.615 7.040 1.845 ;
        RECT  5.345 1.615 5.625 2.095 ;
        RECT  5.345 1.615 5.605 2.120 ;
        RECT  6.755 1.240 7.040 2.690 ;
        RECT  6.755 2.460 8.200 2.690 ;
        RECT  7.860 2.460 8.200 2.800 ;
        RECT  2.905 2.500 3.215 3.115 ;
        RECT  6.635 2.720 6.985 3.295 ;
        RECT  2.905 2.885 4.490 3.115 ;
        RECT  6.755 1.240 6.985 3.295 ;
        RECT  4.260 3.065 6.985 3.295 ;
        RECT  6.295 0.780 7.500 1.010 ;
        RECT  4.885 1.070 5.305 1.385 ;
        RECT  6.295 0.780 6.525 1.385 ;
        RECT  4.885 1.155 6.525 1.385 ;
        RECT  4.885 1.070 5.295 1.390 ;
        RECT  2.640 1.555 3.675 1.785 ;
        RECT  7.270 0.780 7.500 2.020 ;
        RECT  2.640 1.555 2.925 1.895 ;
        RECT  7.270 1.790 8.660 2.020 ;
        RECT  7.990 1.790 8.660 2.130 ;
        RECT  3.445 1.555 3.675 2.655 ;
        RECT  3.445 2.290 3.975 2.655 ;
        RECT  3.445 2.425 5.115 2.655 ;
        RECT  4.885 1.070 5.115 2.655 ;
        RECT  4.905 2.550 5.425 2.835 ;
        RECT  8.430 1.790 8.660 3.240 ;
        RECT  8.430 2.900 8.960 3.240 ;
        RECT  7.730 0.630 10.080 0.950 ;
        RECT  7.730 0.630 8.070 0.970 ;
        RECT  8.510 1.220 8.850 1.560 ;
        RECT  8.510 1.330 9.225 1.560 ;
        RECT  8.995 1.330 9.225 2.635 ;
        RECT  8.995 2.405 10.830 2.635 ;
        RECT  10.130 2.405 10.830 2.745 ;
        RECT  10.130 2.405 10.470 3.375 ;
        RECT  9.290 2.405 9.520 3.820 ;
        RECT  8.340 3.480 9.520 3.820 ;
        RECT  9.460 1.180 11.080 1.410 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  11.070 1.695 11.675 1.980 ;
        RECT  9.460 1.180 9.800 2.010 ;
        RECT  11.070 1.695 11.300 3.205 ;
        RECT  10.770 2.975 11.300 3.205 ;
        RECT  10.770 2.975 11.000 4.180 ;
        RECT  10.600 3.840 11.000 4.180 ;
        RECT  1.220 3.345 2.70 3.575 ;
        RECT  1.635 0.630 3.60 0.860 ;
        RECT  4.260 3.065 5.60 3.295 ;
        RECT  7.730 0.630 9.90 0.950 ;
    END
END DFRRQX1

MACRO DFRRQX0
    CLASS CORE ;
    FOREIGN DFRRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.577  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.315 2.860 11.845 3.350 ;
        RECT  11.615 0.630 11.845 3.350 ;
        RECT  11.180 0.630 11.845 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.245 4.550 2.630 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.500 2.250 10.025 2.815 ;
        END
    END RN
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.200 6.365 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.315 3.810 11.655 5.280 ;
        RECT  9.245 3.910 9.580 5.280 ;
        RECT  6.650 3.630 6.990 5.280 ;
        RECT  4.490 3.910 5.765 5.280 ;
        RECT  0.980 3.520 1.920 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.380 -0.400 10.720 0.950 ;
        RECT  5.710 -0.400 5.995 1.400 ;
        RECT  0.780 -0.400 1.120 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.970 ;
        RECT  0.115 1.740 2.015 1.970 ;
        RECT  1.730 1.740 2.015 2.460 ;
        RECT  0.115 1.360 0.345 3.860 ;
        RECT  0.115 3.520 0.520 3.860 ;
        RECT  2.245 1.285 3.150 1.590 ;
        RECT  0.630 2.200 0.970 3.060 ;
        RECT  0.630 2.720 2.475 3.060 ;
        RECT  2.245 1.285 2.475 4.250 ;
        RECT  2.245 3.910 3.490 4.250 ;
        RECT  1.580 0.825 4.550 1.055 ;
        RECT  1.580 0.825 1.920 1.510 ;
        RECT  4.210 0.825 4.550 1.545 ;
        RECT  5.285 2.160 5.565 2.500 ;
        RECT  6.685 1.230 6.945 3.200 ;
        RECT  2.870 2.840 3.210 3.180 ;
        RECT  5.335 2.860 7.940 3.200 ;
        RECT  2.920 2.840 3.210 3.675 ;
        RECT  5.335 2.160 5.565 3.675 ;
        RECT  2.920 3.445 5.565 3.675 ;
        RECT  6.225 0.765 7.405 0.995 ;
        RECT  4.825 1.230 5.250 1.905 ;
        RECT  4.825 1.675 6.455 1.905 ;
        RECT  6.225 0.765 6.455 1.905 ;
        RECT  3.445 1.775 5.055 2.005 ;
        RECT  7.175 0.765 7.405 2.530 ;
        RECT  2.705 1.835 3.675 2.180 ;
        RECT  7.175 2.170 8.555 2.530 ;
        RECT  3.445 1.775 3.675 3.180 ;
        RECT  4.825 1.230 5.055 3.200 ;
        RECT  3.445 2.860 3.880 3.180 ;
        RECT  4.765 2.860 5.105 3.200 ;
        RECT  8.270 2.170 8.555 3.450 ;
        RECT  7.635 0.630 9.850 0.860 ;
        RECT  7.635 0.630 7.920 0.970 ;
        RECT  9.510 0.630 9.850 0.970 ;
        RECT  8.480 1.170 8.820 1.510 ;
        RECT  8.785 3.125 10.625 3.465 ;
        RECT  8.785 1.280 9.015 3.970 ;
        RECT  7.950 3.680 9.015 3.970 ;
        RECT  11.065 1.360 11.385 1.920 ;
        RECT  9.430 1.690 11.085 2.020 ;
        RECT  10.855 1.690 11.085 4.155 ;
        RECT  10.065 3.925 11.085 4.155 ;
        RECT  10.065 3.925 10.405 4.250 ;
        RECT  1.580 0.825 3.70 1.055 ;
        RECT  5.335 2.860 6.00 3.200 ;
        RECT  2.920 3.445 4.30 3.675 ;
        RECT  7.635 0.630 8.20 0.860 ;
    END
END DFRRQX0

MACRO DFRQX4
    CLASS CORE ;
    FOREIGN DFRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.900 2.250 14.365 2.630 ;
        RECT  13.900 2.250 14.240 3.770 ;
        RECT  11.940 2.250 14.365 2.480 ;
        RECT  13.250 1.130 13.590 2.480 ;
        RECT  12.580 2.250 12.920 3.935 ;
        RECT  11.940 1.095 12.170 2.480 ;
        RECT  11.810 1.095 12.170 1.435 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.550 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.970 -0.400 14.310 1.470 ;
        RECT  12.530 -0.400 12.870 1.470 ;
        RECT  10.310 -0.400 10.650 1.240 ;
        RECT  7.700 -0.400 8.040 1.320 ;
        RECT  5.690 -0.400 6.030 0.950 ;
        RECT  1.580 -0.400 2.400 1.060 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.340 4.170 13.680 5.280 ;
        RECT  11.820 3.910 12.160 5.280 ;
        RECT  10.555 3.540 10.895 5.280 ;
        RECT  8.460 3.850 8.800 5.280 ;
        RECT  6.040 2.910 6.340 5.280 ;
        RECT  1.995 4.060 2.335 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 2.860 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.090 1.190 3.680 1.530 ;
        RECT  1.835 2.325 3.320 2.665 ;
        RECT  3.090 1.190 3.320 3.275 ;
        RECT  3.090 2.935 3.570 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  3.950 2.980 4.290 3.830 ;
        RECT  0.180 3.600 4.290 3.830 ;
        RECT  2.630 0.700 4.140 0.930 ;
        RECT  3.910 0.700 4.140 1.550 ;
        RECT  2.630 0.700 2.860 1.520 ;
        RECT  0.780 1.290 2.860 1.520 ;
        RECT  3.910 1.320 4.495 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.155 1.320 4.495 1.660 ;
        RECT  6.260 0.775 7.470 1.005 ;
        RECT  4.370 0.735 5.295 1.075 ;
        RECT  5.065 0.735 5.295 3.195 ;
        RECT  6.260 0.775 6.490 1.410 ;
        RECT  5.065 1.180 6.490 1.410 ;
        RECT  7.240 0.775 7.470 2.090 ;
        RECT  7.240 1.860 8.950 2.090 ;
        RECT  8.610 1.860 8.950 2.200 ;
        RECT  5.065 1.180 5.350 3.195 ;
        RECT  6.760 1.240 7.010 1.545 ;
        RECT  3.635 1.840 3.975 2.180 ;
        RECT  3.635 1.950 4.835 2.180 ;
        RECT  6.780 1.240 7.010 2.860 ;
        RECT  6.780 2.340 7.830 2.680 ;
        RECT  9.280 1.570 9.565 2.680 ;
        RECT  5.580 2.450 9.565 2.680 ;
        RECT  6.720 2.450 7.060 2.860 ;
        RECT  4.520 1.950 4.835 3.655 ;
        RECT  7.930 3.390 9.550 3.620 ;
        RECT  6.720 2.450 6.950 3.855 ;
        RECT  5.580 2.450 5.810 3.655 ;
        RECT  4.520 3.425 5.810 3.655 ;
        RECT  7.930 3.390 8.160 3.855 ;
        RECT  6.720 3.625 8.160 3.855 ;
        RECT  9.210 3.390 9.550 4.000 ;
        RECT  8.850 0.920 9.190 1.340 ;
        RECT  8.850 1.110 10.025 1.340 ;
        RECT  10.910 2.120 11.250 2.460 ;
        RECT  9.795 2.230 11.250 2.460 ;
        RECT  7.380 2.930 10.025 3.160 ;
        RECT  7.270 3.110 7.610 3.395 ;
        RECT  9.795 1.110 10.025 3.880 ;
        RECT  9.780 2.930 10.025 3.880 ;
        RECT  9.780 3.540 10.120 3.880 ;
        RECT  11.110 0.900 11.450 1.890 ;
        RECT  10.255 1.550 11.450 1.890 ;
        RECT  10.255 1.660 11.710 1.890 ;
        RECT  11.480 1.660 11.710 3.510 ;
        RECT  11.260 2.690 11.710 3.510 ;
        RECT  0.180 3.600 3.70 3.830 ;
        RECT  0.780 1.290 1.70 1.520 ;
        RECT  5.580 2.450 8.60 2.680 ;
        RECT  7.380 2.930 9.50 3.160 ;
    END
END DFRQX4

MACRO DFRQX2
    CLASS CORE ;
    FOREIGN DFRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 1.240 10.600 3.550 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.100 2.100 5.545 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.635 3.770 2.115 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 3.950 11.160 5.280 ;
        RECT  9.500 3.495 9.840 5.280 ;
        RECT  8.295 3.490 8.635 5.280 ;
        RECT  5.910 3.830 6.250 5.280 ;
        RECT  4.770 3.910 5.110 5.280 ;
        RECT  3.510 3.880 3.850 5.280 ;
        RECT  1.680 3.960 2.020 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.820 -0.400 11.160 0.720 ;
        RECT  9.700 -0.400 10.040 0.720 ;
        RECT  8.300 -0.400 8.640 1.060 ;
        RECT  6.650 -0.400 6.990 0.950 ;
        RECT  4.640 -0.400 4.975 0.950 ;
        RECT  3.080 -0.400 3.420 0.840 ;
        RECT  0.700 -0.400 1.040 1.010 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 2.870 ;
        RECT  0.115 2.640 1.455 2.870 ;
        RECT  1.115 2.640 1.455 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  1.270 0.630 2.350 0.950 ;
        RECT  1.270 0.630 1.500 2.410 ;
        RECT  1.270 2.180 1.675 2.410 ;
        RECT  1.625 2.185 1.915 2.415 ;
        RECT  0.575 3.100 0.860 3.440 ;
        RECT  1.685 2.185 1.915 3.625 ;
        RECT  0.575 3.210 1.915 3.440 ;
        RECT  1.685 3.395 2.820 3.625 ;
        RECT  2.480 3.395 2.820 3.735 ;
        RECT  4.460 1.640 5.950 1.870 ;
        RECT  5.665 1.195 5.950 1.870 ;
        RECT  4.460 1.640 4.790 2.180 ;
        RECT  5.775 2.560 6.925 2.900 ;
        RECT  2.145 2.360 2.430 3.165 ;
        RECT  2.145 2.935 3.700 3.165 ;
        RECT  3.470 2.935 3.700 3.410 ;
        RECT  5.530 2.860 6.005 3.410 ;
        RECT  5.775 1.695 6.005 3.410 ;
        RECT  3.470 3.180 6.005 3.410 ;
        RECT  5.205 0.735 6.420 0.965 ;
        RECT  6.190 0.735 6.420 1.555 ;
        RECT  5.205 0.735 5.435 1.410 ;
        RECT  3.880 1.180 5.435 1.410 ;
        RECT  3.880 1.090 4.220 1.430 ;
        RECT  6.190 1.325 7.350 1.555 ;
        RECT  1.730 1.670 2.990 1.955 ;
        RECT  7.120 1.325 7.350 2.190 ;
        RECT  2.760 1.670 2.990 2.705 ;
        RECT  2.760 2.340 3.100 2.705 ;
        RECT  4.000 1.180 4.230 2.950 ;
        RECT  2.760 2.475 4.230 2.705 ;
        RECT  4.000 2.610 4.550 2.950 ;
        RECT  7.265 1.850 7.550 3.310 ;
        RECT  7.475 0.720 8.010 1.060 ;
        RECT  8.920 2.120 9.260 2.460 ;
        RECT  7.780 2.230 9.260 2.460 ;
        RECT  7.780 0.720 8.010 4.005 ;
        RECT  7.065 3.665 8.010 4.005 ;
        RECT  9.000 0.650 9.340 1.180 ;
        RECT  9.000 0.950 9.720 1.180 ;
        RECT  9.490 0.950 9.720 2.960 ;
        RECT  8.240 2.730 9.720 2.960 ;
        RECT  8.240 2.730 9.280 3.070 ;
        RECT  3.470 3.180 5.80 3.410 ;
    END
END DFRQX2

MACRO DFRQX1
    CLASS CORE ;
    FOREIGN DFRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.070 1.030 3.395 2.010 ;
        RECT  2.645 1.030 3.395 1.410 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.695 2.075 5.290 2.360 ;
        RECT  4.535 2.250 4.915 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.662  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.640 2.400 10.585 2.630 ;
        RECT  9.970 2.250 10.585 2.630 ;
        RECT  9.970 1.320 10.200 2.630 ;
        RECT  9.380 1.320 10.200 1.550 ;
        RECT  9.380 3.325 9.870 3.610 ;
        RECT  9.640 2.400 9.870 3.610 ;
        RECT  9.380 0.700 9.720 1.550 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.100 -0.400 10.440 1.090 ;
        RECT  8.575 -0.400 8.915 1.440 ;
        RECT  6.990 -0.400 7.335 0.790 ;
        RECT  4.520 -0.400 4.860 0.925 ;
        RECT  3.060 -0.400 3.400 0.800 ;
        RECT  0.960 -0.400 1.300 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.100 3.330 10.440 5.280 ;
        RECT  8.040 4.145 8.380 5.280 ;
        RECT  5.820 3.810 6.160 5.280 ;
        RECT  4.690 3.525 5.030 5.280 ;
        RECT  3.590 3.810 3.930 5.280 ;
        RECT  1.220 4.170 1.560 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.645 0.520 2.510 ;
        RECT  0.115 2.170 1.020 2.510 ;
        RECT  0.115 0.645 0.345 3.790 ;
        RECT  0.115 3.450 0.760 3.790 ;
        RECT  1.860 0.630 2.200 1.410 ;
        RECT  1.250 1.180 2.200 1.410 ;
        RECT  0.700 2.880 1.480 3.220 ;
        RECT  1.250 1.180 1.480 3.875 ;
        RECT  1.250 3.645 2.530 3.875 ;
        RECT  2.190 3.645 2.530 4.055 ;
        RECT  5.550 1.240 5.835 1.845 ;
        RECT  4.085 1.615 5.835 1.845 ;
        RECT  4.085 1.615 4.365 2.095 ;
        RECT  4.085 1.615 4.345 2.120 ;
        RECT  5.605 1.240 5.835 2.800 ;
        RECT  5.605 2.460 6.870 2.800 ;
        RECT  1.970 2.565 2.310 3.360 ;
        RECT  5.450 2.540 5.810 3.295 ;
        RECT  3.575 3.065 5.810 3.295 ;
        RECT  1.970 3.130 3.755 3.360 ;
        RECT  5.090 0.780 6.295 1.010 ;
        RECT  3.625 1.070 4.100 1.385 ;
        RECT  5.090 0.780 5.320 1.385 ;
        RECT  3.625 1.155 5.320 1.385 ;
        RECT  6.065 0.780 6.295 1.905 ;
        RECT  1.710 1.740 2.050 2.080 ;
        RECT  6.065 1.675 7.130 1.905 ;
        RECT  6.785 1.765 7.505 2.015 ;
        RECT  1.710 1.795 2.840 2.080 ;
        RECT  2.610 1.795 2.840 2.900 ;
        RECT  2.610 2.440 3.855 2.670 ;
        RECT  3.625 1.070 3.855 2.670 ;
        RECT  3.645 2.550 4.230 2.835 ;
        RECT  7.275 1.765 7.505 3.240 ;
        RECT  2.610 2.440 2.980 2.900 ;
        RECT  7.275 2.900 7.630 3.240 ;
        RECT  7.305 1.150 7.645 1.490 ;
        RECT  7.305 1.260 7.965 1.490 ;
        RECT  7.735 1.260 7.965 2.580 ;
        RECT  7.860 2.350 8.940 2.635 ;
        RECT  7.860 2.350 8.090 3.785 ;
        RECT  7.010 3.555 8.090 3.785 ;
        RECT  7.010 3.555 7.350 3.895 ;
        RECT  8.255 1.670 8.595 2.010 ;
        RECT  8.255 1.780 9.720 2.010 ;
        RECT  9.180 1.780 9.720 2.120 ;
        RECT  9.180 1.780 9.410 3.095 ;
        RECT  8.840 2.865 9.410 3.095 ;
        RECT  8.840 2.865 9.150 4.200 ;
        RECT  8.840 3.860 9.180 4.200 ;
        RECT  3.575 3.065 4.20 3.295 ;
    END
END DFRQX1

MACRO DFRQX0
    CLASS CORE ;
    FOREIGN DFRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.493  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.520 2.250 9.955 3.085 ;
        RECT  9.725 0.630 9.955 3.085 ;
        RECT  9.010 0.630 9.955 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 2.220 3.655 2.685 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.000 2.135 5.545 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.445 3.545 9.785 5.280 ;
        RECT  8.040 3.890 8.380 5.280 ;
        RECT  5.300 3.630 5.640 5.280 ;
        RECT  4.420 3.910 4.760 5.280 ;
        RECT  3.490 3.910 3.830 5.280 ;
        RECT  0.780 4.100 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.170 -0.400 8.550 0.970 ;
        RECT  6.510 -0.400 6.795 0.970 ;
        RECT  4.560 -0.400 4.845 0.970 ;
        RECT  3.260 -0.400 3.600 0.970 ;
        RECT  0.780 -0.400 1.120 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.255 0.520 2.395 ;
        RECT  0.115 1.990 1.275 2.395 ;
        RECT  0.115 1.255 0.345 3.700 ;
        RECT  0.115 3.360 0.520 3.700 ;
        RECT  1.505 1.210 2.480 1.505 ;
        RECT  1.505 1.210 1.735 2.775 ;
        RECT  0.575 2.790 1.640 3.020 ;
        RECT  0.575 2.790 0.915 3.130 ;
        RECT  1.410 2.585 1.640 4.230 ;
        RECT  1.410 3.890 2.360 4.230 ;
        RECT  5.535 1.270 5.820 1.905 ;
        RECT  4.345 2.160 4.685 2.500 ;
        RECT  5.775 1.675 6.005 3.200 ;
        RECT  4.455 2.860 6.635 3.200 ;
        RECT  1.870 3.060 2.210 3.400 ;
        RECT  1.980 3.060 2.210 3.660 ;
        RECT  4.455 2.160 4.685 3.660 ;
        RECT  1.980 3.430 4.685 3.660 ;
        RECT  5.075 0.810 6.280 1.040 ;
        RECT  3.885 1.270 4.300 1.610 ;
        RECT  6.050 0.810 6.280 1.445 ;
        RECT  5.075 0.810 5.305 1.610 ;
        RECT  3.885 1.380 5.305 1.610 ;
        RECT  1.965 1.735 4.115 1.965 ;
        RECT  1.965 1.735 2.770 2.080 ;
        RECT  6.235 1.215 6.465 2.460 ;
        RECT  6.235 2.130 6.590 2.460 ;
        RECT  6.235 2.230 7.255 2.460 ;
        RECT  2.540 1.735 2.770 3.180 ;
        RECT  3.885 1.270 4.115 3.200 ;
        RECT  7.010 2.230 7.255 3.425 ;
        RECT  2.540 2.840 2.880 3.180 ;
        RECT  3.820 2.860 4.160 3.200 ;
        RECT  7.010 3.085 7.350 3.425 ;
        RECT  7.310 0.630 7.810 0.970 ;
        RECT  7.580 2.570 8.830 2.910 ;
        RECT  7.580 0.630 7.810 3.970 ;
        RECT  6.700 3.655 7.810 3.970 ;
        RECT  9.010 1.360 9.350 1.700 ;
        RECT  9.010 1.360 9.290 2.130 ;
        RECT  8.060 1.900 9.290 2.130 ;
        RECT  8.060 1.900 8.400 2.240 ;
        RECT  9.060 1.360 9.290 3.370 ;
        RECT  8.555 3.140 9.290 3.370 ;
        RECT  8.555 3.140 8.895 3.480 ;
        RECT  4.455 2.860 5.30 3.200 ;
        RECT  1.980 3.430 3.20 3.660 ;
        RECT  1.965 1.735 3.50 1.965 ;
    END
END DFRQX0

MACRO DFFX4
    CLASS CORE ;
    FOREIGN DFFX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 1.130 16.885 3.770 ;
        RECT  15.170 2.250 16.885 2.630 ;
        RECT  15.170 1.130 15.510 3.935 ;
        RECT  15.050 1.130 15.510 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.078  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.565 2.860 14.890 3.240 ;
        RECT  14.660 1.700 14.890 3.240 ;
        RECT  12.170 1.700 14.890 1.930 ;
        RECT  13.610 1.130 13.950 1.930 ;
        RECT  12.565 2.860 12.945 4.180 ;
        RECT  12.565 2.640 12.930 4.180 ;
        RECT  12.170 1.130 12.510 1.930 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.520 1.640 6.125 2.120 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.770 -0.400 16.110 1.470 ;
        RECT  14.330 -0.400 14.670 1.470 ;
        RECT  12.890 -0.400 13.230 1.470 ;
        RECT  10.310 -0.400 11.090 1.160 ;
        RECT  7.750 -0.400 8.090 1.320 ;
        RECT  5.690 -0.400 6.030 0.950 ;
        RECT  1.580 -0.400 2.400 1.060 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.930 4.170 16.270 5.280 ;
        RECT  14.450 3.555 14.790 5.280 ;
        RECT  13.340 3.870 13.680 5.280 ;
        RECT  11.820 3.910 12.160 5.280 ;
        RECT  10.555 3.540 10.895 5.280 ;
        RECT  8.460 3.850 8.800 5.280 ;
        RECT  6.040 2.910 6.340 5.280 ;
        RECT  0.940 4.060 2.335 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 2.860 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.090 1.190 3.680 1.530 ;
        RECT  1.835 2.325 3.320 2.665 ;
        RECT  3.090 1.190 3.320 3.275 ;
        RECT  3.090 2.935 3.570 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  3.950 2.980 4.290 3.830 ;
        RECT  0.180 3.600 4.290 3.830 ;
        RECT  2.630 0.700 4.140 0.930 ;
        RECT  3.910 0.700 4.140 1.550 ;
        RECT  2.630 0.700 2.860 1.520 ;
        RECT  0.780 1.290 2.860 1.520 ;
        RECT  3.910 1.320 4.495 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.155 1.320 4.495 1.660 ;
        RECT  6.365 0.775 7.520 1.005 ;
        RECT  4.370 0.735 5.295 1.075 ;
        RECT  5.060 0.735 5.295 1.410 ;
        RECT  5.060 1.180 6.600 1.410 ;
        RECT  7.290 0.775 7.520 2.090 ;
        RECT  7.290 1.860 9.000 2.090 ;
        RECT  6.365 0.775 6.600 2.100 ;
        RECT  6.355 1.180 6.600 2.100 ;
        RECT  8.660 1.860 9.000 2.200 ;
        RECT  5.060 0.735 5.290 3.195 ;
        RECT  5.060 2.845 5.350 3.195 ;
        RECT  9.330 1.570 9.620 1.910 ;
        RECT  3.550 1.840 3.860 2.180 ;
        RECT  3.550 1.950 4.830 2.180 ;
        RECT  6.830 2.340 7.830 2.680 ;
        RECT  9.330 1.570 9.560 2.680 ;
        RECT  5.580 2.450 9.560 2.680 ;
        RECT  6.830 1.240 7.060 2.860 ;
        RECT  4.520 1.950 4.830 3.655 ;
        RECT  7.930 3.390 9.550 3.620 ;
        RECT  6.720 2.450 6.950 3.855 ;
        RECT  5.580 2.450 5.810 3.655 ;
        RECT  4.520 3.425 5.810 3.655 ;
        RECT  7.930 3.390 8.160 3.855 ;
        RECT  6.720 3.625 8.160 3.855 ;
        RECT  9.210 3.390 9.550 4.000 ;
        RECT  8.900 0.920 9.240 1.340 ;
        RECT  8.900 1.110 10.080 1.340 ;
        RECT  9.850 1.110 10.080 3.880 ;
        RECT  11.000 1.880 11.340 2.220 ;
        RECT  9.850 1.990 11.340 2.220 ;
        RECT  7.380 2.930 10.120 3.160 ;
        RECT  7.270 3.110 7.610 3.395 ;
        RECT  9.850 1.990 10.120 3.880 ;
        RECT  9.780 2.930 10.120 3.880 ;
        RECT  11.470 0.900 11.810 1.620 ;
        RECT  10.310 1.390 11.810 1.620 ;
        RECT  10.310 1.390 10.650 1.730 ;
        RECT  11.580 2.180 14.430 2.410 ;
        RECT  14.090 2.180 14.430 2.630 ;
        RECT  11.580 0.900 11.810 3.510 ;
        RECT  11.260 2.640 11.810 3.510 ;
        RECT  0.180 3.600 3.10 3.830 ;
        RECT  0.780 1.290 1.40 1.520 ;
        RECT  5.580 2.450 8.80 2.680 ;
        RECT  7.380 2.930 9.40 3.160 ;
        RECT  11.580 2.180 13.40 2.410 ;
    END
END DFFX4

MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.240 11.860 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.200 3.185 11.235 3.415 ;
        RECT  11.005 1.790 11.235 3.415 ;
        RECT  10.200 1.790 11.235 2.020 ;
        RECT  10.200 1.240 10.585 2.020 ;
        RECT  10.200 3.185 10.540 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.635 3.770 2.115 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.470 1.640 4.915 2.030 ;
        RECT  4.470 1.640 4.790 2.180 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  10.960 3.950 12.420 5.280 ;
        RECT  8.295 4.140 9.780 5.280 ;
        RECT  5.910 3.830 6.250 5.280 ;
        RECT  4.770 3.910 5.110 5.280 ;
        RECT  3.510 3.880 3.850 5.280 ;
        RECT  1.680 3.960 2.020 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.960 -0.400 12.420 0.720 ;
        RECT  9.640 -0.400 9.980 0.720 ;
        RECT  8.240 -0.400 8.580 1.130 ;
        RECT  6.650 -0.400 6.990 0.950 ;
        RECT  4.640 -0.400 4.975 0.950 ;
        RECT  3.080 -0.400 3.420 0.840 ;
        RECT  0.700 -0.400 1.040 1.010 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.700 ;
        RECT  0.115 2.640 1.455 2.870 ;
        RECT  1.115 2.640 1.455 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  2.010 0.630 2.350 0.950 ;
        RECT  1.270 0.720 2.350 0.950 ;
        RECT  1.270 0.720 1.500 2.410 ;
        RECT  1.270 2.180 1.675 2.410 ;
        RECT  1.625 2.185 1.915 2.415 ;
        RECT  0.575 3.100 0.860 3.440 ;
        RECT  1.685 2.185 1.915 3.625 ;
        RECT  0.575 3.210 1.915 3.440 ;
        RECT  1.685 3.395 2.820 3.625 ;
        RECT  2.480 3.395 2.820 3.735 ;
        RECT  5.665 1.195 5.950 1.775 ;
        RECT  5.730 1.695 5.960 3.410 ;
        RECT  5.730 2.560 6.925 2.790 ;
        RECT  6.585 2.560 6.925 2.900 ;
        RECT  2.145 2.360 2.430 3.165 ;
        RECT  2.145 2.935 3.700 3.165 ;
        RECT  3.470 2.935 3.700 3.410 ;
        RECT  5.530 2.860 6.005 3.410 ;
        RECT  5.730 2.560 6.005 3.410 ;
        RECT  3.470 3.180 6.005 3.410 ;
        RECT  5.205 0.735 6.420 0.965 ;
        RECT  6.190 0.735 6.420 1.555 ;
        RECT  3.880 1.180 5.435 1.410 ;
        RECT  3.880 1.090 4.220 1.430 ;
        RECT  6.190 1.325 7.290 1.555 ;
        RECT  1.730 1.670 2.990 1.955 ;
        RECT  7.060 1.850 7.400 2.190 ;
        RECT  5.205 0.735 5.435 2.420 ;
        RECT  5.175 1.180 5.435 2.420 ;
        RECT  7.060 1.325 7.290 2.190 ;
        RECT  2.760 1.670 2.990 2.705 ;
        RECT  5.175 2.080 5.500 2.420 ;
        RECT  2.760 2.340 3.100 2.705 ;
        RECT  4.000 1.180 4.230 2.950 ;
        RECT  2.760 2.475 4.230 2.705 ;
        RECT  4.000 2.610 4.550 2.950 ;
        RECT  7.265 1.960 7.550 3.310 ;
        RECT  7.415 0.720 8.010 1.130 ;
        RECT  8.910 2.750 9.250 3.095 ;
        RECT  7.780 2.865 9.250 3.095 ;
        RECT  7.780 0.720 8.010 3.895 ;
        RECT  7.065 3.665 8.010 3.895 ;
        RECT  7.065 3.665 7.405 4.005 ;
        RECT  8.940 0.650 9.280 2.460 ;
        RECT  8.240 2.230 9.710 2.460 ;
        RECT  9.480 2.320 10.775 2.550 ;
        RECT  8.240 2.230 8.580 2.570 ;
        RECT  10.435 2.320 10.775 2.660 ;
        RECT  9.480 2.230 9.710 3.665 ;
        RECT  8.875 3.325 9.710 3.665 ;
        RECT  3.470 3.180 5.30 3.410 ;
    END
END DFFX2

MACRO DFFX1
    CLASS CORE ;
    FOREIGN DFFX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.070 1.670 3.395 2.010 ;
        RECT  3.070 1.180 3.300 2.010 ;
        RECT  2.645 1.180 3.300 1.410 ;
        RECT  2.645 1.030 3.025 1.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.662  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 2.250 10.585 2.630 ;
        RECT  9.640 2.870 10.435 3.100 ;
        RECT  10.205 1.320 10.435 3.100 ;
        RECT  9.490 1.320 10.435 1.550 ;
        RECT  9.380 3.325 9.870 3.610 ;
        RECT  9.640 2.870 9.870 3.610 ;
        RECT  9.490 0.700 9.720 1.550 ;
        RECT  9.380 0.700 9.720 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.820 3.270 11.215 4.180 ;
        RECT  10.820 0.820 11.160 1.160 ;
        RECT  10.820 0.820 11.050 4.180 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.365 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.100 -0.400 10.440 1.090 ;
        RECT  8.575 -0.400 8.915 1.440 ;
        RECT  6.945 -0.400 7.285 0.790 ;
        RECT  4.520 -0.400 4.860 0.925 ;
        RECT  3.060 -0.400 3.400 0.800 ;
        RECT  0.960 -0.400 1.300 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.100 3.330 10.440 5.280 ;
        RECT  8.040 4.145 8.380 5.280 ;
        RECT  5.820 3.810 6.160 5.280 ;
        RECT  4.690 3.525 5.030 5.280 ;
        RECT  3.590 3.810 3.930 5.280 ;
        RECT  1.220 4.170 1.560 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.645 0.520 0.985 ;
        RECT  0.115 2.140 1.020 2.480 ;
        RECT  0.115 0.645 0.345 3.680 ;
        RECT  0.115 3.450 0.760 3.680 ;
        RECT  0.420 3.450 0.760 3.790 ;
        RECT  1.860 0.630 2.200 0.950 ;
        RECT  1.860 0.630 2.090 1.410 ;
        RECT  1.250 1.180 2.090 1.410 ;
        RECT  0.700 2.880 1.480 3.220 ;
        RECT  1.250 1.180 1.480 3.875 ;
        RECT  1.250 3.645 2.530 3.875 ;
        RECT  2.190 3.645 2.530 4.035 ;
        RECT  5.550 1.240 5.835 2.800 ;
        RECT  6.530 2.460 6.870 2.800 ;
        RECT  5.450 2.570 6.870 2.800 ;
        RECT  1.970 2.565 2.310 3.360 ;
        RECT  5.450 2.540 5.810 3.295 ;
        RECT  3.575 3.065 5.810 3.295 ;
        RECT  1.970 3.130 3.755 3.360 ;
        RECT  5.090 0.780 6.295 1.010 ;
        RECT  3.760 1.070 4.100 1.385 ;
        RECT  5.090 0.780 5.320 1.385 ;
        RECT  3.760 1.155 5.320 1.385 ;
        RECT  6.065 0.780 6.295 1.905 ;
        RECT  1.710 1.710 2.050 2.025 ;
        RECT  6.065 1.675 7.130 1.905 ;
        RECT  6.785 1.765 7.505 2.015 ;
        RECT  1.710 1.795 2.840 2.025 ;
        RECT  4.900 1.155 5.290 2.360 ;
        RECT  2.610 1.795 2.840 2.900 ;
        RECT  4.900 1.155 5.130 2.835 ;
        RECT  2.610 2.550 5.130 2.835 ;
        RECT  7.275 1.765 7.505 3.240 ;
        RECT  2.610 2.550 2.980 2.900 ;
        RECT  7.275 2.900 7.630 3.240 ;
        RECT  7.305 1.150 7.645 1.490 ;
        RECT  7.305 1.260 7.965 1.490 ;
        RECT  7.735 1.260 7.965 2.580 ;
        RECT  7.860 2.350 8.940 2.635 ;
        RECT  7.860 2.350 8.090 3.785 ;
        RECT  7.010 3.555 8.090 3.785 ;
        RECT  7.010 3.555 7.350 3.895 ;
        RECT  8.255 1.670 8.595 2.010 ;
        RECT  8.255 1.780 9.720 2.010 ;
        RECT  9.180 1.780 9.720 2.640 ;
        RECT  9.180 2.300 9.870 2.640 ;
        RECT  9.180 1.780 9.410 3.095 ;
        RECT  8.920 2.865 9.410 3.095 ;
        RECT  8.920 2.865 9.150 4.200 ;
        RECT  8.840 3.860 9.180 4.200 ;
        RECT  3.575 3.065 4.20 3.295 ;
        RECT  2.610 2.550 4.50 2.835 ;
    END
END DFFX1

MACRO DFFX0
    CLASS CORE ;
    FOREIGN DFFX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.790 3.710 9.955 3.940 ;
        RECT  9.725 0.630 9.955 3.940 ;
        RECT  9.575 3.470 9.955 3.940 ;
        RECT  9.030 0.630 9.955 0.950 ;
        RECT  8.790 3.710 9.130 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 2.220 3.655 2.685 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.185 1.170 10.585 2.020 ;
        RECT  10.185 3.425 10.530 3.765 ;
        RECT  10.185 1.170 10.415 3.765 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.345 2.160 4.865 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  9.590 4.170 9.930 5.280 ;
        RECT  8.040 3.230 8.325 5.280 ;
        RECT  5.300 3.650 5.640 5.280 ;
        RECT  4.420 3.910 4.760 5.280 ;
        RECT  3.490 3.910 3.830 5.280 ;
        RECT  0.780 4.100 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.190 -0.400 10.530 0.710 ;
        RECT  8.170 -0.400 8.550 0.970 ;
        RECT  6.510 -0.400 6.795 0.970 ;
        RECT  4.560 -0.400 4.845 0.970 ;
        RECT  3.260 -0.400 3.600 0.970 ;
        RECT  0.780 -0.400 1.120 0.965 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.255 0.520 2.410 ;
        RECT  0.115 2.045 1.275 2.410 ;
        RECT  0.115 1.255 0.345 3.700 ;
        RECT  0.115 3.360 0.520 3.700 ;
        RECT  1.505 1.210 2.490 1.505 ;
        RECT  1.505 1.210 1.735 2.795 ;
        RECT  0.575 2.790 1.640 3.020 ;
        RECT  0.575 2.790 0.915 3.130 ;
        RECT  1.410 2.605 1.640 4.230 ;
        RECT  1.410 3.890 2.360 4.230 ;
        RECT  5.555 1.270 5.820 1.905 ;
        RECT  5.665 1.675 5.895 3.200 ;
        RECT  4.455 2.860 6.635 3.200 ;
        RECT  1.870 3.060 2.210 3.400 ;
        RECT  1.980 3.060 2.210 3.660 ;
        RECT  4.455 2.860 4.685 3.660 ;
        RECT  1.980 3.430 4.685 3.660 ;
        RECT  5.075 0.810 6.280 1.040 ;
        RECT  3.885 1.270 4.300 1.610 ;
        RECT  6.050 0.810 6.280 1.445 ;
        RECT  5.075 0.810 5.325 1.610 ;
        RECT  3.885 1.380 5.325 1.610 ;
        RECT  1.965 1.735 4.115 1.965 ;
        RECT  1.965 1.735 2.770 2.100 ;
        RECT  6.235 1.215 6.465 2.480 ;
        RECT  5.095 0.810 5.325 2.575 ;
        RECT  6.235 2.150 6.590 2.480 ;
        RECT  6.235 2.250 7.255 2.480 ;
        RECT  5.095 2.235 5.435 2.575 ;
        RECT  2.540 1.735 2.770 3.180 ;
        RECT  3.885 1.270 4.115 3.200 ;
        RECT  7.010 2.250 7.255 3.470 ;
        RECT  2.540 2.840 2.880 3.180 ;
        RECT  3.820 2.860 4.160 3.200 ;
        RECT  7.010 3.140 7.350 3.470 ;
        RECT  7.330 0.630 7.810 0.970 ;
        RECT  7.580 2.620 8.845 2.960 ;
        RECT  7.580 0.630 7.810 3.990 ;
        RECT  6.535 3.700 7.810 3.990 ;
        RECT  9.030 1.360 9.370 2.180 ;
        RECT  8.080 1.950 9.495 2.180 ;
        RECT  9.075 1.880 9.495 2.220 ;
        RECT  8.080 1.950 8.420 2.290 ;
        RECT  9.075 1.360 9.305 3.480 ;
        RECT  8.790 3.190 9.305 3.480 ;
        RECT  4.455 2.860 5.00 3.200 ;
        RECT  1.980 3.430 3.40 3.660 ;
        RECT  1.965 1.735 3.80 1.965 ;
    END
END DFFX0

MACRO DFFSX4
    CLASS CORE ;
    FOREIGN DFFSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.085  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 1.130 17.460 3.060 ;
        RECT  15.840 2.250 17.460 2.630 ;
        RECT  15.840 2.250 16.180 3.060 ;
        RECT  15.840 1.130 16.070 3.060 ;
        RECT  15.680 1.130 16.070 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.103  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.055 2.890 15.545 3.120 ;
        RECT  15.315 1.700 15.545 3.120 ;
        RECT  12.955 1.700 15.545 1.930 ;
        RECT  13.055 2.890 14.835 3.240 ;
        RECT  14.240 1.130 14.580 1.930 ;
        RECT  13.055 2.860 13.735 3.240 ;
        RECT  13.055 2.860 13.395 4.100 ;
        RECT  12.955 0.630 13.185 1.930 ;
        RECT  12.760 0.630 13.185 0.970 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.255 1.640 11.935 2.020 ;
        RECT  11.255 1.640 11.595 2.220 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.245 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.400 -0.400 16.740 1.470 ;
        RECT  14.960 -0.400 15.300 1.470 ;
        RECT  13.520 -0.400 13.860 1.470 ;
        RECT  10.495 -0.400 11.315 0.880 ;
        RECT  8.115 -0.400 8.455 1.320 ;
        RECT  6.105 -0.400 6.445 0.950 ;
        RECT  1.580 -0.400 2.815 0.710 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.480 3.295 16.820 5.280 ;
        RECT  15.105 3.555 15.445 5.280 ;
        RECT  13.775 3.470 14.115 5.280 ;
        RECT  12.295 4.160 12.635 5.280 ;
        RECT  11.015 3.540 11.355 5.280 ;
        RECT  8.875 3.850 9.215 5.280 ;
        RECT  6.455 2.910 6.755 5.280 ;
        RECT  2.410 3.965 2.750 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 3.275 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.505 1.190 4.095 1.530 ;
        RECT  1.835 2.325 3.735 2.665 ;
        RECT  3.505 1.190 3.735 3.275 ;
        RECT  3.505 2.935 3.985 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.650 3.735 ;
        RECT  4.365 2.980 4.650 3.735 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  3.045 0.700 4.555 0.930 ;
        RECT  4.325 0.700 4.555 1.550 ;
        RECT  3.045 0.700 3.275 1.520 ;
        RECT  0.780 1.290 3.275 1.520 ;
        RECT  4.325 1.320 4.910 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.570 1.320 4.910 1.660 ;
        RECT  6.675 0.775 7.885 1.005 ;
        RECT  4.785 0.735 5.645 1.075 ;
        RECT  5.335 0.735 5.645 1.410 ;
        RECT  5.335 1.180 6.905 1.410 ;
        RECT  6.675 0.775 6.905 2.100 ;
        RECT  6.625 1.180 6.905 2.100 ;
        RECT  7.655 0.775 7.885 2.090 ;
        RECT  7.655 1.860 9.365 2.090 ;
        RECT  6.625 1.760 6.910 2.100 ;
        RECT  9.025 1.860 9.365 2.200 ;
        RECT  5.335 0.735 5.565 2.375 ;
        RECT  5.340 2.275 5.570 3.195 ;
        RECT  5.340 2.855 5.765 3.195 ;
        RECT  7.170 1.240 7.425 1.555 ;
        RECT  9.695 1.570 10.020 1.910 ;
        RECT  7.195 1.240 7.425 2.860 ;
        RECT  7.195 2.340 8.245 2.680 ;
        RECT  3.965 1.840 4.275 2.705 ;
        RECT  9.695 1.570 9.925 2.680 ;
        RECT  5.995 2.450 9.925 2.680 ;
        RECT  3.965 2.475 5.110 2.705 ;
        RECT  7.135 2.450 7.475 2.860 ;
        RECT  4.880 2.475 5.110 3.655 ;
        RECT  8.345 3.390 9.965 3.620 ;
        RECT  7.135 2.450 7.365 3.855 ;
        RECT  5.995 2.450 6.225 3.655 ;
        RECT  4.880 3.425 6.225 3.655 ;
        RECT  8.345 3.390 8.575 3.855 ;
        RECT  7.135 3.625 8.575 3.855 ;
        RECT  9.625 3.390 9.965 4.000 ;
        RECT  9.265 0.920 9.605 1.340 ;
        RECT  9.265 1.110 10.480 1.340 ;
        RECT  10.250 1.110 10.480 3.880 ;
        RECT  11.925 2.370 12.265 2.710 ;
        RECT  10.250 2.480 12.265 2.710 ;
        RECT  7.795 2.930 10.535 3.160 ;
        RECT  7.685 3.110 8.025 3.395 ;
        RECT  10.250 2.480 10.535 3.880 ;
        RECT  10.195 2.930 10.535 3.880 ;
        RECT  10.710 1.140 12.505 1.370 ;
        RECT  10.710 1.140 10.995 1.480 ;
        RECT  12.165 1.140 12.505 1.620 ;
        RECT  12.495 2.310 15.085 2.540 ;
        RECT  14.745 2.310 15.085 2.650 ;
        RECT  12.495 1.390 12.725 3.170 ;
        RECT  11.735 2.940 12.725 3.170 ;
        RECT  11.735 2.940 12.075 3.760 ;
        RECT  2.030 3.505 3.40 3.735 ;
        RECT  0.180 3.600 1.90 3.830 ;
        RECT  0.780 1.290 2.40 1.520 ;
        RECT  5.995 2.450 8.90 2.680 ;
        RECT  10.250 2.480 11.30 2.710 ;
        RECT  7.795 2.930 9.20 3.160 ;
        RECT  12.495 2.310 14.80 2.540 ;
    END
END DFFSX4

MACRO DFFSX2
    CLASS CORE ;
    FOREIGN DFFSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.090 1.640 5.545 2.140 ;
        END
    END CN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 1.240 13.120 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.899  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.460 2.860 12.495 3.090 ;
        RECT  12.265 1.180 12.495 3.090 ;
        RECT  11.460 1.180 12.495 1.410 ;
        RECT  11.460 0.840 11.845 1.410 ;
        RECT  11.460 2.860 11.800 4.180 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.800 2.250 10.585 2.705 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 1.630 4.400 2.110 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.220 3.950 13.680 5.280 ;
        RECT  10.715 3.940 11.055 5.280 ;
        RECT  9.235 3.865 9.575 5.280 ;
        RECT  6.940 3.470 7.280 5.280 ;
        RECT  5.640 3.525 5.980 5.280 ;
        RECT  4.340 3.525 4.680 5.280 ;
        RECT  1.700 3.910 2.550 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.220 -0.400 13.680 0.720 ;
        RECT  10.740 -0.400 11.080 1.060 ;
        RECT  9.205 -0.400 9.545 1.090 ;
        RECT  7.280 -0.400 7.620 0.890 ;
        RECT  5.270 -0.400 5.610 0.950 ;
        RECT  3.640 -0.400 3.980 0.825 ;
        RECT  1.130 -0.400 1.470 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.700 ;
        RECT  0.115 2.585 2.040 2.815 ;
        RECT  1.730 2.585 2.040 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  1.700 1.035 2.780 1.325 ;
        RECT  1.700 1.035 1.930 2.355 ;
        RECT  1.700 2.125 2.500 2.355 ;
        RECT  0.575 3.100 0.915 3.440 ;
        RECT  2.270 2.125 2.500 3.575 ;
        RECT  0.575 3.210 2.500 3.440 ;
        RECT  2.270 3.345 3.350 3.575 ;
        RECT  3.010 3.345 3.350 3.685 ;
        RECT  6.300 1.240 6.590 1.580 ;
        RECT  6.360 1.240 6.590 3.295 ;
        RECT  6.360 2.280 8.035 2.510 ;
        RECT  7.695 2.280 8.035 2.605 ;
        RECT  2.730 2.310 3.060 2.650 ;
        RECT  2.830 2.310 3.060 3.115 ;
        RECT  2.830 2.885 4.330 3.115 ;
        RECT  6.360 2.280 6.740 3.295 ;
        RECT  4.100 3.065 6.740 3.295 ;
        RECT  5.840 0.780 7.050 1.010 ;
        RECT  4.510 1.070 4.850 1.410 ;
        RECT  4.510 1.180 6.070 1.410 ;
        RECT  2.160 1.555 2.500 1.895 ;
        RECT  6.820 0.780 7.050 1.900 ;
        RECT  5.840 0.780 6.070 2.100 ;
        RECT  5.790 1.180 6.070 2.100 ;
        RECT  2.160 1.665 3.620 1.895 ;
        RECT  6.820 1.670 7.545 1.900 ;
        RECT  7.205 1.780 8.495 2.010 ;
        RECT  5.790 1.760 6.130 2.100 ;
        RECT  3.390 1.665 3.620 2.655 ;
        RECT  3.390 2.290 3.730 2.655 ;
        RECT  4.630 1.180 4.860 2.835 ;
        RECT  3.390 2.425 4.860 2.655 ;
        RECT  4.630 2.550 5.220 2.835 ;
        RECT  8.265 1.780 8.495 3.065 ;
        RECT  7.635 2.835 8.495 3.065 ;
        RECT  7.635 2.835 7.865 4.040 ;
        RECT  7.635 3.810 8.795 4.040 ;
        RECT  8.485 3.805 8.795 4.100 ;
        RECT  8.455 3.810 8.795 4.100 ;
        RECT  8.175 0.630 8.955 0.950 ;
        RECT  8.725 2.965 10.720 3.250 ;
        RECT  8.725 0.630 8.955 3.525 ;
        RECT  8.095 3.295 8.955 3.525 ;
        RECT  8.095 3.295 8.435 3.580 ;
        RECT  10.540 1.560 10.880 2.020 ;
        RECT  9.185 1.790 11.180 2.020 ;
        RECT  10.950 2.120 12.035 2.460 ;
        RECT  9.185 1.790 9.470 2.700 ;
        RECT  10.950 1.790 11.180 3.710 ;
        RECT  9.965 3.480 11.180 3.710 ;
        RECT  9.965 3.480 10.305 4.070 ;
        RECT  4.100 3.065 5.60 3.295 ;
    END
END DFFSX2

MACRO DFFSX1
    CLASS CORE ;
    FOREIGN DFFSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.630 2.100 ;
        END
    END CN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.475 2.085 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.640 10.585 2.305 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 2.250 12.475 2.630 ;
        RECT  11.530 2.870 12.325 3.100 ;
        RECT  12.095 1.235 12.325 3.100 ;
        RECT  11.380 1.235 12.325 1.465 ;
        RECT  11.270 3.665 11.760 4.005 ;
        RECT  11.530 2.870 11.760 4.005 ;
        RECT  11.380 0.700 11.610 1.465 ;
        RECT  11.270 0.700 11.610 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 0.820 13.105 4.180 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.990 -0.400 12.330 1.005 ;
        RECT  10.015 -0.400 10.355 0.880 ;
        RECT  7.725 -0.400 8.065 0.820 ;
        RECT  5.665 -0.400 6.005 0.950 ;
        RECT  4.165 -0.400 4.475 1.410 ;
        RECT  1.340 -0.400 1.680 1.565 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  11.990 3.330 12.330 5.280 ;
        RECT  10.570 4.005 10.910 5.280 ;
        RECT  9.210 3.910 9.550 5.280 ;
        RECT  7.110 3.320 7.450 5.280 ;
        RECT  5.810 3.525 6.150 5.280 ;
        RECT  4.510 3.525 4.850 5.280 ;
        RECT  1.670 3.820 2.015 5.280 ;
        RECT  0.180 3.870 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.025 ;
        RECT  0.170 1.795 1.815 2.025 ;
        RECT  1.475 1.795 1.815 2.135 ;
        RECT  0.780 1.795 1.120 3.085 ;
        RECT  2.045 1.175 2.940 1.515 ;
        RECT  0.260 3.235 0.600 3.575 ;
        RECT  2.045 1.175 2.275 3.575 ;
        RECT  0.260 3.345 3.450 3.575 ;
        RECT  3.110 3.345 3.450 3.665 ;
        RECT  6.695 1.240 7.035 1.580 ;
        RECT  6.695 2.310 8.125 2.540 ;
        RECT  7.785 2.310 8.125 2.650 ;
        RECT  6.695 1.240 6.925 2.880 ;
        RECT  2.625 2.500 2.965 3.115 ;
        RECT  6.560 2.540 6.790 3.295 ;
        RECT  2.625 2.885 4.425 3.115 ;
        RECT  4.195 3.065 6.790 3.295 ;
        RECT  6.235 0.780 7.495 1.010 ;
        RECT  4.705 1.070 5.245 1.410 ;
        RECT  4.705 1.180 6.465 1.410 ;
        RECT  7.265 0.780 7.495 1.870 ;
        RECT  7.265 1.640 8.325 1.870 ;
        RECT  7.985 1.695 8.690 1.980 ;
        RECT  2.505 1.745 3.675 2.085 ;
        RECT  6.235 0.780 6.465 2.100 ;
        RECT  6.075 1.760 6.465 2.100 ;
        RECT  3.445 1.745 3.675 2.655 ;
        RECT  3.445 2.315 3.900 2.655 ;
        RECT  4.705 1.070 4.935 2.835 ;
        RECT  3.445 2.425 4.935 2.655 ;
        RECT  8.460 1.695 8.690 3.080 ;
        RECT  4.705 2.550 5.350 2.835 ;
        RECT  8.460 2.740 8.800 3.080 ;
        RECT  8.505 1.110 9.225 1.450 ;
        RECT  8.995 1.110 9.225 2.460 ;
        RECT  9.035 2.635 10.830 2.975 ;
        RECT  9.035 2.230 9.265 3.550 ;
        RECT  8.380 3.320 9.265 3.550 ;
        RECT  8.380 3.320 8.720 4.250 ;
        RECT  9.455 1.180 11.080 1.410 ;
        RECT  9.455 1.180 9.795 1.720 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  11.070 1.695 11.570 2.500 ;
        RECT  11.070 2.160 11.725 2.500 ;
        RECT  11.070 1.695 11.300 3.435 ;
        RECT  9.970 3.205 11.300 3.435 ;
        RECT  9.970 3.205 10.310 3.605 ;
        RECT  0.260 3.345 2.30 3.575 ;
        RECT  4.195 3.065 5.20 3.295 ;
    END
END DFFSX1

MACRO DFFSX0
    CLASS CORE ;
    FOREIGN DFFSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.975 2.250 5.495 2.630 ;
        RECT  4.975 2.165 5.315 2.630 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.645 2.715 11.215 3.240 ;
        RECT  10.985 0.630 11.215 3.240 ;
        RECT  10.070 0.630 11.215 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.760 2.220 4.285 2.685 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.360 2.210 9.955 2.630 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.502  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.445 1.170 11.845 3.765 ;
        END
    END QN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  10.645 3.515 10.985 5.280 ;
        RECT  8.690 3.635 9.030 5.280 ;
        RECT  6.095 3.630 6.435 5.280 ;
        RECT  5.050 3.910 5.390 5.280 ;
        RECT  4.120 3.910 4.460 5.280 ;
        RECT  1.470 3.360 1.810 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  11.450 -0.400 11.790 0.710 ;
        RECT  8.970 -0.400 9.315 0.970 ;
        RECT  7.140 -0.400 7.425 0.970 ;
        RECT  5.190 -0.400 5.475 0.970 ;
        RECT  3.890 -0.400 4.230 0.990 ;
        RECT  1.300 -0.400 1.640 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.270 0.630 0.610 1.930 ;
        RECT  0.115 1.700 1.905 1.930 ;
        RECT  1.620 1.700 1.905 2.080 ;
        RECT  0.115 1.700 0.345 3.060 ;
        RECT  0.115 2.770 1.080 3.060 ;
        RECT  0.740 2.770 1.080 3.700 ;
        RECT  2.690 1.165 3.030 1.505 ;
        RECT  2.135 1.275 3.030 1.505 ;
        RECT  0.575 2.200 0.860 2.540 ;
        RECT  2.135 1.275 2.365 2.540 ;
        RECT  0.575 2.310 2.365 2.540 ;
        RECT  2.040 2.310 2.270 4.140 ;
        RECT  2.040 3.910 3.120 4.140 ;
        RECT  2.780 3.910 3.120 4.250 ;
        RECT  6.165 1.270 6.450 3.200 ;
        RECT  2.500 2.840 2.840 3.180 ;
        RECT  5.635 2.860 7.385 3.200 ;
        RECT  2.610 2.840 2.840 3.675 ;
        RECT  5.635 2.860 5.865 3.675 ;
        RECT  2.610 3.445 5.865 3.675 ;
        RECT  5.705 0.810 6.910 1.040 ;
        RECT  4.515 1.270 5.935 1.500 ;
        RECT  4.515 1.270 4.930 1.610 ;
        RECT  2.595 1.735 4.745 1.965 ;
        RECT  2.595 1.735 3.400 2.080 ;
        RECT  5.705 0.810 5.935 2.130 ;
        RECT  6.680 0.810 6.910 2.350 ;
        RECT  6.865 2.120 8.000 2.460 ;
        RECT  3.170 1.735 3.400 3.180 ;
        RECT  4.515 1.270 4.745 3.200 ;
        RECT  3.170 2.840 3.510 3.180 ;
        RECT  4.450 2.860 4.790 3.200 ;
        RECT  7.715 2.120 8.000 3.425 ;
        RECT  7.940 0.630 8.460 0.970 ;
        RECT  8.230 2.880 9.955 3.110 ;
        RECT  9.640 2.880 9.955 3.220 ;
        RECT  8.230 0.630 8.460 3.970 ;
        RECT  7.435 3.655 8.460 3.970 ;
        RECT  8.690 1.690 10.410 1.920 ;
        RECT  10.070 1.310 10.410 1.920 ;
        RECT  8.690 1.690 9.030 2.105 ;
        RECT  10.185 1.830 10.755 2.170 ;
        RECT  10.185 1.830 10.415 3.970 ;
        RECT  9.475 3.630 10.415 3.970 ;
        RECT  2.610 3.445 4.50 3.675 ;
        RECT  2.595 1.735 3.00 1.965 ;
    END
END DFFSX0

MACRO DFFSQX4
    CLASS CORE ;
    FOREIGN DFFSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.600 1.130 14.940 4.130 ;
        RECT  13.280 2.250 14.940 2.630 ;
        RECT  13.280 0.790 13.620 2.630 ;
        RECT  13.160 2.890 13.510 4.100 ;
        RECT  13.280 0.790 13.510 4.100 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.110 1.640 11.845 2.020 ;
        RECT  11.110 1.640 11.450 2.090 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.245 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.120 0.400 ;
        RECT  14.040 -0.400 14.380 0.720 ;
        RECT  12.520 -0.400 12.860 0.710 ;
        RECT  10.825 -0.400 11.165 0.910 ;
        RECT  8.060 -0.400 8.345 1.320 ;
        RECT  6.105 -0.400 6.445 0.950 ;
        RECT  1.580 -0.400 2.815 0.710 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.120 5.280 ;
        RECT  13.880 2.890 14.220 5.280 ;
        RECT  12.400 4.160 12.740 5.280 ;
        RECT  11.015 3.540 11.355 5.280 ;
        RECT  8.875 3.850 9.215 5.280 ;
        RECT  6.455 2.910 6.755 5.280 ;
        RECT  2.410 3.965 2.750 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 3.275 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.505 1.190 4.095 1.530 ;
        RECT  1.835 2.325 3.735 2.665 ;
        RECT  3.505 1.190 3.735 3.275 ;
        RECT  3.505 2.935 3.985 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.650 3.735 ;
        RECT  4.365 2.980 4.650 3.735 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  3.045 0.700 4.555 0.930 ;
        RECT  4.325 0.700 4.555 1.550 ;
        RECT  3.045 0.700 3.275 1.520 ;
        RECT  0.780 1.290 3.275 1.520 ;
        RECT  4.325 1.320 4.910 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.570 1.320 4.910 1.660 ;
        RECT  6.675 0.775 7.830 1.005 ;
        RECT  4.785 0.735 5.645 1.075 ;
        RECT  5.335 0.735 5.645 1.410 ;
        RECT  5.335 1.180 6.905 1.410 ;
        RECT  7.600 0.775 7.830 1.910 ;
        RECT  6.675 0.775 6.905 2.100 ;
        RECT  6.625 1.180 6.905 2.100 ;
        RECT  7.600 1.680 9.255 1.910 ;
        RECT  8.915 1.680 9.255 2.020 ;
        RECT  6.625 1.760 6.910 2.100 ;
        RECT  5.335 0.735 5.565 2.375 ;
        RECT  5.340 2.275 5.570 3.195 ;
        RECT  5.340 2.855 5.765 3.195 ;
        RECT  7.135 1.240 7.370 1.580 ;
        RECT  7.140 1.240 7.370 2.860 ;
        RECT  7.140 2.340 7.995 2.680 ;
        RECT  3.965 1.840 4.275 2.705 ;
        RECT  9.585 1.520 9.870 2.680 ;
        RECT  5.995 2.450 9.870 2.680 ;
        RECT  3.965 2.475 5.110 2.705 ;
        RECT  7.135 2.450 7.475 2.860 ;
        RECT  4.880 2.475 5.110 3.655 ;
        RECT  8.345 3.390 9.965 3.620 ;
        RECT  7.135 2.450 7.365 3.855 ;
        RECT  5.995 2.450 6.225 3.655 ;
        RECT  4.880 3.425 6.225 3.655 ;
        RECT  8.345 3.390 8.575 3.855 ;
        RECT  7.135 3.625 8.575 3.855 ;
        RECT  9.625 3.390 9.965 4.000 ;
        RECT  9.155 0.920 9.495 1.290 ;
        RECT  9.155 1.060 10.330 1.290 ;
        RECT  11.925 2.370 12.265 2.710 ;
        RECT  10.100 2.480 12.265 2.710 ;
        RECT  7.795 2.930 10.425 3.160 ;
        RECT  10.100 1.060 10.330 3.160 ;
        RECT  7.685 3.110 8.025 3.395 ;
        RECT  10.195 2.480 10.425 3.880 ;
        RECT  10.195 3.540 10.535 3.880 ;
        RECT  10.560 1.140 12.360 1.370 ;
        RECT  10.560 1.140 10.845 1.480 ;
        RECT  12.020 1.250 12.725 1.480 ;
        RECT  12.495 1.250 12.725 3.170 ;
        RECT  11.735 2.940 12.725 3.170 ;
        RECT  11.735 2.940 12.075 3.760 ;
        RECT  2.030 3.505 3.40 3.735 ;
        RECT  0.180 3.600 1.60 3.830 ;
        RECT  0.780 1.290 2.50 1.520 ;
        RECT  5.995 2.450 8.10 2.680 ;
        RECT  10.100 2.480 11.40 2.710 ;
        RECT  7.795 2.930 9.60 3.160 ;
    END
END DFFSQX4

MACRO DFFSQX2
    CLASS CORE ;
    FOREIGN DFFSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.180 11.860 3.550 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.800 2.250 10.585 2.735 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 1.630 4.400 2.110 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.090 1.640 5.545 2.140 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  10.960 3.995 12.420 5.280 ;
        RECT  9.425 3.425 9.765 5.280 ;
        RECT  6.940 3.470 7.280 5.280 ;
        RECT  5.640 3.525 5.980 5.280 ;
        RECT  4.340 3.525 4.680 5.280 ;
        RECT  1.700 3.910 2.550 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.960 -0.400 12.420 0.720 ;
        RECT  9.205 -0.400 9.545 1.090 ;
        RECT  7.280 -0.400 7.620 0.890 ;
        RECT  5.270 -0.400 5.610 0.950 ;
        RECT  3.640 -0.400 3.980 0.825 ;
        RECT  1.130 -0.400 1.470 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.700 ;
        RECT  0.115 2.585 2.040 2.815 ;
        RECT  1.730 2.585 2.040 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  1.700 1.035 2.780 1.325 ;
        RECT  1.700 1.035 1.930 2.355 ;
        RECT  1.700 2.125 2.500 2.355 ;
        RECT  0.575 3.100 0.915 3.440 ;
        RECT  2.270 2.125 2.500 3.575 ;
        RECT  0.575 3.210 2.500 3.440 ;
        RECT  2.270 3.345 3.350 3.575 ;
        RECT  3.010 3.345 3.350 3.685 ;
        RECT  6.300 1.240 6.590 1.580 ;
        RECT  6.360 1.240 6.590 3.295 ;
        RECT  6.360 2.280 8.035 2.510 ;
        RECT  7.695 2.280 8.035 2.605 ;
        RECT  2.730 2.310 3.060 2.650 ;
        RECT  2.830 2.310 3.060 3.115 ;
        RECT  2.830 2.885 4.330 3.115 ;
        RECT  6.360 2.280 6.740 3.295 ;
        RECT  4.100 3.065 6.740 3.295 ;
        RECT  5.840 0.780 7.050 1.010 ;
        RECT  4.510 1.070 4.850 1.410 ;
        RECT  4.510 1.180 6.070 1.410 ;
        RECT  2.160 1.555 2.500 1.895 ;
        RECT  6.820 0.780 7.050 1.900 ;
        RECT  5.840 0.780 6.070 2.100 ;
        RECT  5.790 1.180 6.070 2.100 ;
        RECT  2.160 1.665 3.620 1.895 ;
        RECT  6.820 1.670 7.545 1.900 ;
        RECT  7.205 1.780 8.495 2.010 ;
        RECT  5.790 1.760 6.130 2.100 ;
        RECT  3.390 1.665 3.620 2.655 ;
        RECT  3.390 2.290 3.730 2.655 ;
        RECT  4.630 1.180 4.860 2.835 ;
        RECT  3.390 2.425 4.860 2.655 ;
        RECT  4.630 2.550 5.220 2.835 ;
        RECT  8.265 1.780 8.495 3.065 ;
        RECT  7.635 2.835 8.495 3.065 ;
        RECT  7.635 2.835 7.865 4.040 ;
        RECT  7.635 3.810 8.795 4.040 ;
        RECT  8.455 3.810 8.795 4.100 ;
        RECT  8.175 0.630 8.955 0.950 ;
        RECT  8.725 2.965 10.775 3.195 ;
        RECT  10.435 2.965 10.775 3.305 ;
        RECT  8.725 0.630 8.955 3.580 ;
        RECT  8.095 3.295 8.955 3.580 ;
        RECT  10.235 0.680 10.575 2.020 ;
        RECT  9.185 1.790 11.235 2.020 ;
        RECT  9.185 1.790 9.470 2.700 ;
        RECT  11.005 1.790 11.235 3.765 ;
        RECT  10.200 3.535 11.235 3.765 ;
        RECT  10.200 3.535 10.540 4.070 ;
        RECT  4.100 3.065 5.40 3.295 ;
        RECT  8.725 2.965 9.80 3.195 ;
        RECT  9.185 1.790 10.40 2.020 ;
    END
END DFFSQX2

MACRO DFFSQX1
    CLASS CORE ;
    FOREIGN DFFSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.475 2.085 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.110 1.640 10.585 2.305 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.530 2.400 12.475 2.630 ;
        RECT  11.800 2.250 12.475 2.630 ;
        RECT  11.800 1.235 12.030 2.630 ;
        RECT  11.380 1.235 12.030 1.465 ;
        RECT  11.270 3.665 11.760 4.005 ;
        RECT  11.530 2.400 11.760 4.005 ;
        RECT  11.380 0.700 11.610 1.465 ;
        RECT  11.270 0.700 11.610 1.040 ;
        END
    END Q
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.630 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  11.990 -0.400 12.330 1.005 ;
        RECT  10.015 -0.400 10.355 0.880 ;
        RECT  7.725 -0.400 8.065 0.790 ;
        RECT  5.665 -0.400 6.005 0.950 ;
        RECT  4.165 -0.400 4.475 1.410 ;
        RECT  1.340 -0.400 1.680 1.565 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.990 3.330 12.330 5.280 ;
        RECT  10.570 4.005 10.910 5.280 ;
        RECT  9.210 3.910 9.550 5.280 ;
        RECT  7.110 3.320 7.450 5.280 ;
        RECT  5.810 3.525 6.150 5.280 ;
        RECT  4.510 3.525 4.850 5.280 ;
        RECT  1.670 3.820 2.015 5.280 ;
        RECT  0.180 3.870 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.025 ;
        RECT  0.170 1.795 1.815 2.025 ;
        RECT  1.475 1.795 1.815 2.135 ;
        RECT  0.780 1.795 1.120 3.085 ;
        RECT  2.045 1.175 2.940 1.515 ;
        RECT  0.260 3.235 0.600 3.575 ;
        RECT  2.045 1.175 2.275 3.575 ;
        RECT  0.260 3.345 3.450 3.575 ;
        RECT  3.110 3.345 3.450 3.665 ;
        RECT  6.695 1.240 7.035 1.580 ;
        RECT  6.695 2.310 8.125 2.540 ;
        RECT  7.785 2.310 8.125 2.650 ;
        RECT  6.695 1.240 6.925 2.880 ;
        RECT  2.645 2.500 2.985 3.115 ;
        RECT  6.560 2.540 6.790 3.295 ;
        RECT  2.645 2.885 4.425 3.115 ;
        RECT  4.195 3.065 6.790 3.295 ;
        RECT  6.235 0.780 7.495 1.010 ;
        RECT  4.705 1.070 5.245 1.410 ;
        RECT  4.705 1.180 6.465 1.410 ;
        RECT  7.265 0.780 7.495 1.870 ;
        RECT  7.265 1.640 8.325 1.870 ;
        RECT  7.985 1.695 8.690 1.980 ;
        RECT  2.505 1.745 3.675 2.085 ;
        RECT  6.235 0.780 6.465 2.100 ;
        RECT  6.075 1.760 6.465 2.100 ;
        RECT  3.445 1.745 3.675 2.655 ;
        RECT  3.445 2.315 3.900 2.655 ;
        RECT  4.705 1.070 4.935 2.835 ;
        RECT  3.445 2.425 4.935 2.655 ;
        RECT  8.460 1.695 8.690 3.080 ;
        RECT  4.705 2.550 5.350 2.835 ;
        RECT  8.460 2.740 8.800 3.080 ;
        RECT  8.505 1.110 9.225 1.450 ;
        RECT  8.995 1.110 9.225 2.460 ;
        RECT  9.035 2.635 10.830 2.865 ;
        RECT  10.490 2.635 10.830 2.975 ;
        RECT  9.035 2.230 9.265 3.550 ;
        RECT  8.380 3.320 9.265 3.550 ;
        RECT  8.380 3.320 8.720 4.250 ;
        RECT  9.455 1.180 11.080 1.410 ;
        RECT  9.455 1.180 9.795 1.720 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  11.070 1.695 11.570 1.980 ;
        RECT  11.070 1.695 11.300 3.435 ;
        RECT  9.970 3.205 11.300 3.435 ;
        RECT  9.970 3.205 10.310 3.605 ;
        RECT  0.260 3.345 2.40 3.575 ;
        RECT  4.195 3.065 5.30 3.295 ;
    END
END DFFSQX1

MACRO DFFSQX0
    CLASS CORE ;
    FOREIGN DFFSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.975 2.250 5.495 2.630 ;
        RECT  4.975 2.165 5.315 2.630 ;
        END
    END CN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.542  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.670 2.715 11.215 3.240 ;
        RECT  10.985 0.630 11.215 3.240 ;
        RECT  10.200 0.630 11.215 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.760 2.220 4.285 2.685 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.360 2.210 9.955 2.630 ;
        END
    END SN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.670 3.515 11.010 5.280 ;
        RECT  8.690 3.635 9.030 5.280 ;
        RECT  6.095 3.630 6.435 5.280 ;
        RECT  5.050 3.910 5.390 5.280 ;
        RECT  4.120 3.910 4.460 5.280 ;
        RECT  1.470 3.360 1.810 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  8.970 -0.400 9.315 1.420 ;
        RECT  7.140 -0.400 7.425 0.970 ;
        RECT  5.190 -0.400 5.475 0.970 ;
        RECT  3.890 -0.400 4.230 0.990 ;
        RECT  1.300 -0.400 1.640 1.470 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.270 0.630 0.610 1.930 ;
        RECT  0.115 1.700 1.905 1.930 ;
        RECT  1.620 1.700 1.905 2.080 ;
        RECT  0.115 1.700 0.345 3.060 ;
        RECT  0.115 2.770 1.080 3.060 ;
        RECT  0.740 2.770 1.080 3.700 ;
        RECT  2.690 1.165 3.030 1.505 ;
        RECT  2.135 1.275 3.030 1.505 ;
        RECT  0.575 2.200 0.860 2.540 ;
        RECT  2.135 1.275 2.365 2.540 ;
        RECT  0.575 2.310 2.365 2.540 ;
        RECT  2.040 2.310 2.270 4.140 ;
        RECT  2.040 3.910 3.120 4.140 ;
        RECT  2.780 3.910 3.120 4.250 ;
        RECT  6.165 1.270 6.450 3.200 ;
        RECT  2.500 2.840 2.840 3.180 ;
        RECT  5.635 2.860 7.385 3.200 ;
        RECT  2.610 2.840 2.840 3.675 ;
        RECT  5.635 2.860 5.865 3.675 ;
        RECT  2.610 3.445 5.865 3.675 ;
        RECT  5.705 0.810 6.910 1.040 ;
        RECT  4.515 1.270 5.935 1.500 ;
        RECT  4.515 1.270 4.930 1.610 ;
        RECT  2.595 1.735 4.745 1.965 ;
        RECT  2.595 1.735 3.400 2.080 ;
        RECT  5.705 0.810 5.935 2.130 ;
        RECT  6.680 0.810 6.910 2.460 ;
        RECT  6.680 2.170 8.000 2.460 ;
        RECT  3.170 1.735 3.400 3.180 ;
        RECT  4.515 1.270 4.745 3.200 ;
        RECT  3.170 2.840 3.510 3.180 ;
        RECT  4.450 2.860 4.790 3.200 ;
        RECT  7.715 2.170 8.000 3.425 ;
        RECT  7.940 0.630 8.460 0.970 ;
        RECT  8.230 2.880 9.955 3.110 ;
        RECT  9.640 2.880 9.955 3.220 ;
        RECT  8.230 0.630 8.460 3.970 ;
        RECT  7.435 3.655 8.460 3.970 ;
        RECT  10.200 1.310 10.540 1.650 ;
        RECT  8.690 1.690 10.440 1.920 ;
        RECT  8.690 1.690 9.030 2.105 ;
        RECT  10.185 1.690 10.440 3.970 ;
        RECT  10.200 1.310 10.440 3.970 ;
        RECT  9.510 3.630 10.440 3.970 ;
        RECT  2.610 3.445 4.20 3.675 ;
        RECT  2.595 1.735 3.80 1.965 ;
    END
END DFFSQX0

MACRO DFFRX4
    CLASS CORE ;
    FOREIGN DFFRX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.931  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.380 1.130 18.775 3.260 ;
        RECT  17.180 2.250 18.775 2.630 ;
        RECT  17.180 2.250 17.560 3.240 ;
        RECT  17.180 1.130 17.410 3.240 ;
        RECT  16.940 1.130 17.410 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.078  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 2.880 16.950 3.220 ;
        RECT  16.720 1.700 16.950 3.220 ;
        RECT  14.170 1.700 16.950 1.930 ;
        RECT  15.500 1.130 15.840 1.930 ;
        RECT  14.615 2.640 14.995 4.180 ;
        RECT  14.170 1.130 14.400 1.930 ;
        RECT  14.060 1.130 14.400 1.470 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.290 1.640 13.105 2.020 ;
        RECT  12.290 1.640 12.630 2.190 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.760 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.670 1.660 7.435 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  17.660 -0.400 18.000 1.470 ;
        RECT  16.220 -0.400 16.560 1.470 ;
        RECT  14.780 -0.400 15.120 1.470 ;
        RECT  12.800 -0.400 13.140 0.710 ;
        RECT  7.230 -0.400 7.515 0.970 ;
        RECT  1.750 -0.400 3.225 0.655 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  17.800 3.625 18.130 5.280 ;
        RECT  16.640 3.580 16.980 5.280 ;
        RECT  15.390 3.870 15.730 5.280 ;
        RECT  13.870 4.110 14.210 5.280 ;
        RECT  11.490 3.760 12.950 5.280 ;
        RECT  9.315 4.170 9.655 5.280 ;
        RECT  6.825 3.925 7.165 5.280 ;
        RECT  2.410 3.985 3.245 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.805 1.920 2.090 ;
        RECT  1.375 1.860 3.420 2.090 ;
        RECT  3.190 1.860 3.420 2.800 ;
        RECT  3.190 2.460 3.530 2.800 ;
        RECT  1.375 1.805 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.780 1.345 3.935 1.575 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  2.325 1.345 3.935 1.630 ;
        RECT  3.645 1.345 3.935 1.695 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.525 5.200 3.755 ;
        RECT  4.860 3.010 5.200 3.755 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  4.165 1.160 5.210 1.500 ;
        RECT  1.835 2.325 2.580 2.665 ;
        RECT  4.165 1.160 4.395 3.295 ;
        RECT  2.240 2.325 2.580 3.295 ;
        RECT  4.140 2.955 4.480 3.295 ;
        RECT  2.240 3.065 4.480 3.295 ;
        RECT  0.180 0.640 0.520 1.015 ;
        RECT  3.520 0.700 5.670 0.930 ;
        RECT  0.180 0.785 1.520 1.015 ;
        RECT  1.290 0.885 3.750 1.115 ;
        RECT  5.440 0.700 5.670 1.660 ;
        RECT  5.440 1.320 5.980 1.660 ;
        RECT  7.745 0.775 8.895 1.005 ;
        RECT  5.900 0.735 6.770 1.090 ;
        RECT  6.210 0.735 6.770 1.430 ;
        RECT  6.210 1.200 7.975 1.430 ;
        RECT  8.665 0.775 8.895 2.090 ;
        RECT  8.665 1.860 10.330 2.090 ;
        RECT  9.990 1.860 10.330 2.200 ;
        RECT  7.745 0.775 7.975 2.225 ;
        RECT  7.665 1.200 7.975 2.225 ;
        RECT  6.210 0.735 6.440 3.235 ;
        RECT  6.050 2.895 6.440 3.235 ;
        RECT  4.625 1.890 5.810 2.120 ;
        RECT  8.205 1.240 8.435 2.805 ;
        RECT  8.205 2.340 8.685 2.805 ;
        RECT  8.205 2.520 10.945 2.805 ;
        RECT  10.660 1.670 10.945 2.805 ;
        RECT  7.585 2.575 10.945 2.805 ;
        RECT  7.585 2.575 7.925 2.915 ;
        RECT  5.470 1.890 5.810 3.695 ;
        RECT  5.470 3.465 7.815 3.695 ;
        RECT  7.585 2.575 7.815 3.940 ;
        RECT  7.585 3.710 10.170 3.940 ;
        RECT  9.940 3.710 10.170 4.250 ;
        RECT  9.940 3.965 10.280 4.250 ;
        RECT  9.125 0.630 12.340 0.860 ;
        RECT  11.530 0.630 12.340 0.950 ;
        RECT  9.125 0.630 9.420 1.500 ;
        RECT  10.230 1.100 10.570 1.440 ;
        RECT  10.230 1.210 11.405 1.440 ;
        RECT  11.175 1.210 11.405 3.395 ;
        RECT  13.140 2.310 13.480 2.650 ;
        RECT  11.175 2.420 13.480 2.650 ;
        RECT  12.050 2.420 12.390 3.150 ;
        RECT  11.175 2.420 11.460 3.395 ;
        RECT  8.125 3.165 11.460 3.395 ;
        RECT  8.125 3.165 8.465 3.480 ;
        RECT  10.485 3.165 10.800 3.860 ;
        RECT  10.510 3.165 10.800 3.890 ;
        RECT  11.635 1.180 13.700 1.410 ;
        RECT  13.360 1.110 13.700 1.905 ;
        RECT  11.635 1.180 11.975 1.675 ;
        RECT  13.360 1.675 13.940 1.905 ;
        RECT  13.710 2.180 16.480 2.410 ;
        RECT  16.140 2.180 16.480 2.650 ;
        RECT  13.710 1.675 13.940 3.110 ;
        RECT  13.310 2.880 13.940 3.110 ;
        RECT  13.310 2.880 13.650 3.700 ;
        RECT  1.375 1.860 2.80 2.090 ;
        RECT  0.780 1.345 2.80 1.575 ;
        RECT  2.030 3.525 4.30 3.755 ;
        RECT  0.180 3.600 1.70 3.830 ;
        RECT  2.240 3.065 3.30 3.295 ;
        RECT  3.520 0.700 4.70 0.930 ;
        RECT  1.290 0.885 2.10 1.115 ;
        RECT  8.205 2.520 9.30 2.805 ;
        RECT  7.585 2.575 9.20 2.805 ;
        RECT  5.470 3.465 6.80 3.695 ;
        RECT  7.585 3.710 9.60 3.940 ;
        RECT  9.125 0.630 11.60 0.860 ;
        RECT  11.175 2.420 12.90 2.650 ;
        RECT  8.125 3.165 10.80 3.395 ;
        RECT  11.635 1.180 12.20 1.410 ;
        RECT  13.710 2.180 15.80 2.410 ;
    END
END DFFRX4

MACRO DFFRX2
    CLASS CORE ;
    FOREIGN DFFRX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 1.240 13.750 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.090 2.860 13.105 3.090 ;
        RECT  12.875 0.950 13.105 3.090 ;
        RECT  12.090 0.950 13.105 1.180 ;
        RECT  12.090 2.860 12.475 4.180 ;
        RECT  12.090 0.820 12.430 1.180 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.080 1.940 10.585 2.630 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.400 1.640 4.915 2.120 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 1.640 5.585 2.140 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  12.850 3.950 14.310 5.280 ;
        RECT  11.370 3.785 11.710 5.280 ;
        RECT  9.620 3.860 9.960 5.280 ;
        RECT  7.200 3.660 7.540 5.280 ;
        RECT  5.900 3.525 6.240 5.280 ;
        RECT  4.600 3.525 4.940 5.280 ;
        RECT  1.470 3.805 2.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  12.850 -0.400 14.310 0.720 ;
        RECT  11.330 -0.400 11.670 0.720 ;
        RECT  10.430 -0.400 10.770 0.710 ;
        RECT  5.390 -0.400 5.730 0.950 ;
        RECT  0.780 -0.400 1.120 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.360 0.520 2.510 ;
        RECT  0.115 2.280 1.905 2.510 ;
        RECT  1.620 2.280 1.905 2.620 ;
        RECT  0.115 2.280 0.345 4.070 ;
        RECT  0.115 3.730 0.620 4.070 ;
        RECT  2.700 1.305 3.040 1.645 ;
        RECT  2.135 1.415 3.040 1.645 ;
        RECT  0.575 2.850 2.365 3.190 ;
        RECT  2.135 1.415 2.365 3.575 ;
        RECT  2.135 3.345 3.630 3.575 ;
        RECT  3.290 3.345 3.630 3.685 ;
        RECT  1.580 0.630 4.240 0.950 ;
        RECT  1.580 0.630 1.920 1.090 ;
        RECT  6.425 1.240 6.850 1.580 ;
        RECT  6.620 1.240 6.850 3.295 ;
        RECT  7.920 2.360 8.260 2.700 ;
        RECT  6.620 2.470 8.260 2.700 ;
        RECT  3.010 2.505 3.350 3.115 ;
        RECT  3.010 2.885 4.910 3.115 ;
        RECT  6.620 2.470 7.000 3.295 ;
        RECT  4.680 3.065 7.000 3.295 ;
        RECT  5.965 0.780 7.310 1.010 ;
        RECT  4.630 1.070 5.070 1.410 ;
        RECT  3.680 1.180 6.195 1.410 ;
        RECT  7.080 0.780 7.310 1.980 ;
        RECT  7.080 1.750 7.660 1.980 ;
        RECT  5.965 0.780 6.195 2.365 ;
        RECT  7.320 1.860 8.740 2.090 ;
        RECT  2.595 1.880 3.910 2.220 ;
        RECT  3.680 1.180 3.910 2.655 ;
        RECT  5.965 2.020 6.390 2.365 ;
        RECT  3.680 2.315 4.020 2.655 ;
        RECT  3.680 2.425 5.480 2.655 ;
        RECT  8.510 1.860 8.740 3.130 ;
        RECT  5.140 2.425 5.480 2.835 ;
        RECT  8.510 2.790 9.010 3.130 ;
        RECT  7.540 0.630 10.010 0.970 ;
        RECT  9.670 0.630 10.010 1.040 ;
        RECT  8.440 1.210 9.200 1.550 ;
        RECT  8.970 1.210 9.200 2.200 ;
        RECT  8.970 1.970 9.550 2.200 ;
        RECT  9.320 2.860 11.135 3.090 ;
        RECT  10.795 2.750 11.135 3.095 ;
        RECT  10.180 2.860 11.135 3.095 ;
        RECT  10.180 2.860 10.520 3.200 ;
        RECT  9.320 1.970 9.550 3.630 ;
        RECT  8.385 3.400 9.550 3.630 ;
        RECT  8.385 3.400 8.725 3.825 ;
        RECT  9.430 1.400 11.670 1.630 ;
        RECT  9.430 1.400 9.770 1.740 ;
        RECT  11.330 1.400 11.670 1.980 ;
        RECT  11.440 2.120 12.645 2.460 ;
        RECT  11.440 1.400 11.670 3.555 ;
        RECT  10.760 3.325 11.670 3.555 ;
        RECT  10.760 3.325 10.990 4.125 ;
        RECT  10.650 3.785 10.990 4.125 ;
        RECT  1.580 0.630 3.30 0.950 ;
        RECT  4.680 3.065 6.70 3.295 ;
        RECT  3.680 1.180 5.30 1.410 ;
        RECT  7.540 0.630 9.70 0.970 ;
        RECT  9.430 1.400 10.90 1.630 ;
    END
END DFFRX2

MACRO DFFRX1
    CLASS CORE ;
    FOREIGN DFFRX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.630 2.100 ;
        END
    END CN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.655 2.025 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.050 1.640 10.610 2.085 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.678  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 2.250 12.475 2.630 ;
        RECT  11.530 2.870 12.325 3.100 ;
        RECT  12.095 1.235 12.325 3.100 ;
        RECT  11.380 1.235 12.325 1.465 ;
        RECT  11.270 3.435 11.760 3.720 ;
        RECT  11.530 2.870 11.760 3.720 ;
        RECT  11.380 0.700 11.610 1.465 ;
        RECT  11.270 0.700 11.610 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.710 0.820 13.105 4.180 ;
        END
    END QN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.990 -0.400 12.330 1.005 ;
        RECT  10.470 -0.400 10.810 0.950 ;
        RECT  5.725 -0.400 6.065 0.930 ;
        RECT  0.915 -0.400 1.255 1.395 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  11.990 3.330 12.330 5.280 ;
        RECT  9.800 3.850 10.140 5.280 ;
        RECT  7.185 3.480 7.525 5.280 ;
        RECT  5.885 3.525 6.225 5.280 ;
        RECT  4.585 3.525 4.925 5.280 ;
        RECT  1.940 3.840 2.280 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.215 0.645 0.555 2.350 ;
        RECT  0.115 2.120 1.950 2.350 ;
        RECT  1.665 2.120 1.950 2.460 ;
        RECT  0.115 2.120 0.345 3.790 ;
        RECT  0.115 3.450 0.760 3.790 ;
        RECT  2.180 1.090 3.205 1.325 ;
        RECT  0.575 2.855 1.555 3.195 ;
        RECT  1.220 2.855 1.555 4.180 ;
        RECT  2.180 1.090 2.410 3.575 ;
        RECT  1.220 3.345 3.525 3.575 ;
        RECT  3.185 3.345 3.525 3.665 ;
        RECT  1.220 3.345 1.560 4.180 ;
        RECT  1.635 0.630 4.605 0.860 ;
        RECT  4.265 0.630 4.605 1.280 ;
        RECT  1.635 0.630 1.950 1.450 ;
        RECT  6.755 1.240 7.040 2.690 ;
        RECT  6.755 2.460 8.200 2.690 ;
        RECT  7.860 2.460 8.200 2.800 ;
        RECT  2.905 2.290 3.215 3.115 ;
        RECT  6.635 2.720 6.985 3.295 ;
        RECT  2.905 2.885 4.490 3.115 ;
        RECT  6.755 1.240 6.985 3.295 ;
        RECT  4.260 3.065 6.985 3.295 ;
        RECT  6.295 0.780 7.500 1.010 ;
        RECT  4.960 1.070 5.305 1.390 ;
        RECT  6.295 0.780 6.525 1.385 ;
        RECT  4.960 1.160 6.365 1.390 ;
        RECT  2.640 1.555 3.675 1.785 ;
        RECT  7.270 0.780 7.500 2.020 ;
        RECT  2.640 1.555 2.925 1.895 ;
        RECT  7.270 1.790 8.660 2.020 ;
        RECT  7.990 1.790 8.660 2.130 ;
        RECT  6.100 1.900 6.490 2.240 ;
        RECT  3.445 1.555 3.675 2.655 ;
        RECT  3.445 2.290 3.975 2.655 ;
        RECT  6.100 1.160 6.365 2.655 ;
        RECT  3.445 2.425 6.365 2.655 ;
        RECT  5.080 2.425 5.425 2.835 ;
        RECT  8.430 1.790 8.660 3.240 ;
        RECT  8.430 2.900 8.960 3.240 ;
        RECT  7.730 0.630 10.010 0.860 ;
        RECT  9.670 0.630 10.010 0.950 ;
        RECT  7.730 0.630 8.070 0.970 ;
        RECT  8.510 1.220 9.225 1.560 ;
        RECT  8.995 1.220 9.225 2.635 ;
        RECT  8.995 2.405 10.840 2.635 ;
        RECT  10.130 2.405 10.840 2.745 ;
        RECT  10.130 2.405 10.470 3.385 ;
        RECT  9.290 2.405 9.520 3.820 ;
        RECT  8.340 3.480 9.520 3.820 ;
        RECT  9.460 1.180 11.080 1.410 ;
        RECT  9.460 1.180 9.800 2.025 ;
        RECT  10.850 1.695 11.610 2.175 ;
        RECT  10.850 1.180 11.080 2.175 ;
        RECT  11.070 2.160 11.865 2.500 ;
        RECT  11.070 1.695 11.300 3.205 ;
        RECT  10.770 2.975 11.300 3.205 ;
        RECT  10.770 2.975 11.000 4.190 ;
        RECT  10.600 3.850 11.000 4.190 ;
        RECT  1.220 3.345 2.70 3.575 ;
        RECT  1.635 0.630 3.80 0.860 ;
        RECT  4.260 3.065 5.30 3.295 ;
        RECT  3.445 2.425 5.20 2.655 ;
        RECT  7.730 0.630 9.80 0.860 ;
    END
END DFFRX1

MACRO DFFRX0
    CLASS CORE ;
    FOREIGN DFFRX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.577  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.315 2.860 11.875 3.350 ;
        RECT  11.645 0.630 11.875 3.350 ;
        RECT  11.180 0.630 11.875 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.245 4.525 2.630 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.500 2.250 10.025 2.815 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.441  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.105 1.170 12.475 4.150 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.215 2.200 5.680 2.645 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.315 3.810 11.655 5.280 ;
        RECT  9.245 3.910 9.580 5.280 ;
        RECT  6.650 3.630 6.990 5.280 ;
        RECT  4.490 3.910 5.765 5.280 ;
        RECT  0.980 3.520 1.920 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.105 -0.400 12.420 0.710 ;
        RECT  10.380 -0.400 10.720 0.950 ;
        RECT  5.710 -0.400 5.995 1.400 ;
        RECT  0.780 -0.400 1.120 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.970 ;
        RECT  0.115 1.740 2.015 1.970 ;
        RECT  1.730 1.740 2.015 2.460 ;
        RECT  0.115 1.360 0.345 3.860 ;
        RECT  0.115 3.520 0.520 3.860 ;
        RECT  2.245 1.285 3.150 1.590 ;
        RECT  0.630 2.200 0.970 3.060 ;
        RECT  0.630 2.720 2.475 3.060 ;
        RECT  2.245 1.285 2.475 4.140 ;
        RECT  2.245 3.910 3.490 4.140 ;
        RECT  3.110 3.910 3.490 4.250 ;
        RECT  1.580 0.825 4.550 1.055 ;
        RECT  1.580 0.825 1.920 1.510 ;
        RECT  4.210 0.825 4.550 1.545 ;
        RECT  6.685 1.230 6.945 3.200 ;
        RECT  2.870 2.840 3.210 3.180 ;
        RECT  6.225 2.860 7.940 3.200 ;
        RECT  5.335 2.900 7.940 3.200 ;
        RECT  2.920 2.840 3.210 3.675 ;
        RECT  5.335 2.900 5.565 3.675 ;
        RECT  2.920 3.445 5.565 3.675 ;
        RECT  6.225 0.765 7.405 0.995 ;
        RECT  4.825 1.230 5.250 1.950 ;
        RECT  4.825 1.720 6.455 1.950 ;
        RECT  6.225 0.765 6.455 1.950 ;
        RECT  3.445 1.775 4.985 2.005 ;
        RECT  7.175 0.765 7.405 2.530 ;
        RECT  2.705 1.835 3.675 2.180 ;
        RECT  7.175 2.170 8.555 2.530 ;
        RECT  5.990 1.720 6.330 2.575 ;
        RECT  3.445 1.775 3.675 3.180 ;
        RECT  4.755 1.775 4.985 3.200 ;
        RECT  3.445 2.860 3.880 3.180 ;
        RECT  4.755 2.860 5.105 3.200 ;
        RECT  8.270 2.170 8.555 3.450 ;
        RECT  7.635 0.630 9.850 0.860 ;
        RECT  7.635 0.630 7.920 0.970 ;
        RECT  9.510 0.630 9.850 0.970 ;
        RECT  8.480 1.170 8.820 1.510 ;
        RECT  8.785 3.125 10.625 3.465 ;
        RECT  8.785 1.280 9.015 3.970 ;
        RECT  7.950 3.680 9.015 3.970 ;
        RECT  9.430 1.690 11.415 1.920 ;
        RECT  9.430 1.690 9.770 2.020 ;
        RECT  11.065 1.360 11.415 2.220 ;
        RECT  10.855 1.690 11.085 4.155 ;
        RECT  10.065 3.925 11.085 4.155 ;
        RECT  10.065 3.925 10.405 4.250 ;
        RECT  1.580 0.825 3.60 1.055 ;
        RECT  5.335 2.900 6.40 3.200 ;
        RECT  2.920 3.445 4.90 3.675 ;
        RECT  7.635 0.630 8.40 0.860 ;
    END
END DFFRX0

MACRO DFFRSX4
    CLASS CORE ;
    FOREIGN DFFRSX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.105  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 1.130 19.980 3.295 ;
        RECT  18.345 2.250 19.980 2.630 ;
        RECT  18.345 2.250 18.685 3.295 ;
        RECT  18.345 1.130 18.575 3.295 ;
        RECT  18.200 1.130 18.575 1.470 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.135  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.635 3.010 18.065 3.240 ;
        RECT  17.835 1.700 18.065 3.240 ;
        RECT  15.580 1.700 18.065 1.930 ;
        RECT  17.075 3.010 17.415 3.350 ;
        RECT  16.760 1.130 17.100 1.930 ;
        RECT  15.635 2.860 16.255 3.240 ;
        RECT  15.635 2.860 15.975 4.030 ;
        RECT  15.580 1.130 15.810 1.930 ;
        RECT  15.320 1.130 15.810 1.470 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.905 1.640 14.365 2.525 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.725 2.250 13.485 2.630 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.600 1.660 8.065 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.920 -0.400 19.260 1.470 ;
        RECT  17.480 -0.400 17.820 1.470 ;
        RECT  16.040 -0.400 16.380 1.470 ;
        RECT  13.430 -0.400 13.770 0.950 ;
        RECT  7.830 -0.400 8.115 0.970 ;
        RECT  2.255 -0.400 3.825 0.665 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  19.000 3.530 19.340 5.280 ;
        RECT  17.705 3.685 18.045 5.280 ;
        RECT  16.355 3.470 16.695 5.280 ;
        RECT  14.875 4.060 15.215 5.280 ;
        RECT  12.435 3.910 13.895 5.280 ;
        RECT  10.135 3.965 10.475 5.280 ;
        RECT  7.715 2.910 8.015 5.280 ;
        RECT  2.410 3.965 3.845 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.765 1.815 2.105 2.095 ;
        RECT  1.375 1.860 4.020 2.095 ;
        RECT  3.790 1.860 4.020 2.800 ;
        RECT  3.790 2.460 4.130 2.800 ;
        RECT  1.375 1.860 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.965 1.355 4.535 1.585 ;
        RECT  0.965 1.290 1.305 1.630 ;
        RECT  2.925 1.355 4.535 1.630 ;
        RECT  4.245 1.355 4.535 1.695 ;
        RECT  5.475 1.160 5.810 1.500 ;
        RECT  4.765 1.270 5.810 1.500 ;
        RECT  1.835 2.325 3.180 2.665 ;
        RECT  2.840 2.325 3.180 3.275 ;
        RECT  4.765 1.270 4.995 3.540 ;
        RECT  2.840 3.045 4.995 3.275 ;
        RECT  4.735 3.200 5.080 3.540 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.415 3.735 ;
        RECT  4.185 3.505 4.415 4.000 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  5.500 2.980 5.840 4.000 ;
        RECT  4.185 3.770 5.840 4.000 ;
        RECT  0.365 0.640 0.705 1.015 ;
        RECT  4.120 0.630 6.270 0.860 ;
        RECT  0.365 0.785 2.025 1.015 ;
        RECT  4.120 0.630 4.350 1.125 ;
        RECT  1.795 0.895 4.350 1.125 ;
        RECT  6.040 0.630 6.270 1.660 ;
        RECT  6.040 1.320 6.625 1.660 ;
        RECT  8.345 0.775 9.495 1.005 ;
        RECT  6.500 0.735 7.370 1.090 ;
        RECT  7.140 1.200 8.575 1.430 ;
        RECT  9.265 0.775 9.495 2.090 ;
        RECT  9.265 1.860 10.930 2.090 ;
        RECT  8.345 0.775 8.575 2.100 ;
        RECT  8.295 1.200 8.575 2.100 ;
        RECT  7.140 0.735 7.370 2.150 ;
        RECT  6.795 1.920 7.370 2.150 ;
        RECT  10.590 1.860 10.930 2.200 ;
        RECT  6.795 1.920 7.025 3.195 ;
        RECT  6.685 2.855 7.025 3.195 ;
        RECT  5.225 1.820 5.565 2.120 ;
        RECT  11.260 1.670 11.600 2.010 ;
        RECT  5.225 1.890 6.455 2.120 ;
        RECT  8.805 1.240 9.035 2.680 ;
        RECT  8.805 2.340 9.505 2.680 ;
        RECT  11.260 1.670 11.490 2.680 ;
        RECT  7.255 2.450 11.490 2.680 ;
        RECT  8.395 2.450 8.735 2.860 ;
        RECT  6.225 1.890 6.455 3.655 ;
        RECT  8.395 2.450 8.625 3.855 ;
        RECT  7.255 2.450 7.485 3.655 ;
        RECT  6.225 3.425 7.485 3.655 ;
        RECT  9.605 3.505 11.225 3.735 ;
        RECT  8.395 3.625 9.835 3.855 ;
        RECT  10.885 3.505 11.225 4.100 ;
        RECT  9.725 0.630 12.965 0.860 ;
        RECT  1.375 1.860 3.60 2.095 ;
        RECT  0.965 1.355 3.50 1.585 ;
        RECT  2.840 3.045 3.30 3.275 ;
        RECT  2.030 3.505 3.40 3.735 ;
        RECT  0.180 3.600 1.60 3.830 ;
        RECT  4.120 0.630 5.50 0.860 ;
        RECT  1.795 0.895 3.20 1.125 ;
        RECT  7.255 2.450 10.60 2.680 ;
        RECT  9.725 0.630 11.40 0.860 ;
        RECT  12.155 0.630 12.965 0.950 ;
        RECT  9.725 0.630 10.020 1.500 ;
        RECT  10.830 1.100 11.170 1.440 ;
        RECT  10.830 1.210 12.060 1.440 ;
        RECT  11.830 1.210 12.060 3.275 ;
        RECT  12.995 2.860 14.890 3.090 ;
        RECT  14.595 2.270 14.890 3.090 ;
        RECT  8.945 3.045 13.335 3.275 ;
        RECT  8.945 3.045 9.285 3.395 ;
        RECT  11.455 3.045 11.745 3.980 ;
        RECT  12.290 1.180 14.960 1.410 ;
        RECT  14.620 1.080 14.960 1.420 ;
        RECT  12.290 1.180 12.630 1.730 ;
        RECT  14.730 1.080 14.960 2.040 ;
        RECT  14.730 1.810 15.350 2.040 ;
        RECT  15.120 2.250 17.605 2.480 ;
        RECT  17.265 2.250 17.605 2.590 ;
        RECT  15.120 1.810 15.350 3.550 ;
        RECT  14.315 3.320 15.350 3.550 ;
        RECT  14.315 3.320 14.655 3.660 ;
    END
END DFFRSX4

MACRO DFFRSX2
    CLASS CORE ;
    FOREIGN DFFRSX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  14.615 1.240 15.010 3.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.350 2.860 14.365 3.090 ;
        RECT  14.135 0.950 14.365 3.090 ;
        RECT  13.350 0.950 14.365 1.180 ;
        RECT  13.350 2.860 13.735 4.180 ;
        RECT  13.350 0.820 13.690 1.180 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.790 1.920 11.215 2.630 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.445 1.640 11.915 2.160 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.820 1.640 5.105 2.100 ;
        RECT  4.535 1.640 5.105 2.020 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.290 2.100 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  14.110 3.950 15.570 5.280 ;
        RECT  12.630 3.785 12.970 5.280 ;
        RECT  11.190 3.730 11.530 5.280 ;
        RECT  10.200 3.860 10.540 5.280 ;
        RECT  7.730 3.480 8.070 5.280 ;
        RECT  6.430 3.525 6.770 5.280 ;
        RECT  5.130 3.525 5.470 5.280 ;
        RECT  1.500 3.805 2.900 5.280 ;
        RECT  0.180 3.780 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  14.110 -0.400 15.570 0.720 ;
        RECT  12.590 -0.400 12.930 0.720 ;
        RECT  11.155 -0.400 11.495 0.710 ;
        RECT  6.060 -0.400 6.400 0.950 ;
        RECT  1.210 -0.400 1.550 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.360 0.520 2.070 ;
        RECT  0.130 1.840 2.405 2.070 ;
        RECT  2.120 1.840 2.405 2.490 ;
        RECT  0.130 1.360 0.360 3.160 ;
        RECT  0.130 2.870 1.080 3.160 ;
        RECT  2.635 1.090 3.540 1.325 ;
        RECT  0.590 2.300 0.930 2.640 ;
        RECT  0.590 2.410 1.630 2.640 ;
        RECT  1.400 2.410 1.630 3.190 ;
        RECT  1.400 2.850 2.865 3.190 ;
        RECT  2.635 1.090 2.865 3.575 ;
        RECT  2.635 3.345 3.930 3.575 ;
        RECT  3.590 3.345 3.930 3.820 ;
        RECT  1.970 0.630 4.940 0.860 ;
        RECT  4.600 0.630 4.940 1.410 ;
        RECT  1.970 0.630 2.310 1.530 ;
        RECT  7.090 1.240 7.380 1.580 ;
        RECT  7.150 1.240 7.380 3.295 ;
        RECT  7.150 2.320 8.865 2.550 ;
        RECT  8.525 2.320 8.865 2.660 ;
        RECT  3.510 2.310 3.845 3.115 ;
        RECT  3.510 2.885 5.020 3.115 ;
        RECT  7.150 2.320 7.530 3.295 ;
        RECT  4.790 3.065 7.530 3.295 ;
        RECT  6.630 0.780 7.840 1.010 ;
        RECT  5.300 1.070 5.640 1.410 ;
        RECT  5.300 1.180 6.860 1.410 ;
        RECT  7.610 0.780 7.840 1.940 ;
        RECT  6.630 0.780 6.860 2.100 ;
        RECT  6.580 1.180 6.860 2.100 ;
        RECT  3.095 1.555 4.305 1.895 ;
        RECT  7.610 1.710 8.385 1.940 ;
        RECT  8.045 1.820 9.325 2.050 ;
        RECT  6.580 1.760 6.920 2.100 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 4.520 2.655 ;
        RECT  5.335 1.070 5.565 2.835 ;
        RECT  4.075 2.425 5.565 2.655 ;
        RECT  9.095 1.820 9.325 3.090 ;
        RECT  5.335 2.550 6.010 2.835 ;
        RECT  9.095 2.750 9.590 3.090 ;
        RECT  8.070 0.630 10.735 0.860 ;
        RECT  8.070 0.630 8.355 0.970 ;
        RECT  10.395 0.630 10.735 1.015 ;
        RECT  10.395 0.630 10.725 1.030 ;
        RECT  9.165 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  9.820 2.860 12.650 3.090 ;
        RECT  12.310 2.750 12.650 3.095 ;
        RECT  10.760 2.860 12.650 3.095 ;
        RECT  10.760 2.860 11.100 3.200 ;
        RECT  9.820 1.970 10.050 3.550 ;
        RECT  8.970 3.320 10.050 3.550 ;
        RECT  8.970 3.320 9.310 3.660 ;
        RECT  10.900 1.180 12.930 1.410 ;
        RECT  10.115 1.400 11.130 1.630 ;
        RECT  10.115 1.400 10.455 1.740 ;
        RECT  12.590 1.180 12.930 1.980 ;
        RECT  12.890 2.120 13.905 2.460 ;
        RECT  12.890 1.695 13.120 3.555 ;
        RECT  11.910 3.325 13.120 3.555 ;
        RECT  11.910 3.325 12.250 4.070 ;
        RECT  0.130 1.840 1.80 2.070 ;
        RECT  1.970 0.630 3.80 0.860 ;
        RECT  4.790 3.065 6.70 3.295 ;
        RECT  8.070 0.630 9.00 0.860 ;
        RECT  9.820 2.860 11.60 3.090 ;
        RECT  10.900 1.180 11.50 1.410 ;
    END
END DFFRSX2

MACRO DFFRSX1
    CLASS CORE ;
    FOREIGN DFFRSX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.105 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.640 11.845 2.305 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.835 2.045 11.215 2.630 ;
        RECT  10.520 2.045 11.215 2.385 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.710  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 2.250 13.735 2.630 ;
        RECT  12.790 2.870 13.585 3.100 ;
        RECT  13.355 1.235 13.585 3.100 ;
        RECT  12.640 1.235 13.585 1.465 ;
        RECT  12.530 3.630 13.020 3.915 ;
        RECT  12.790 2.870 13.020 3.915 ;
        RECT  12.640 0.700 12.870 1.465 ;
        RECT  12.530 0.700 12.870 1.040 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.792  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.970 3.270 14.365 4.180 ;
        RECT  13.970 0.820 14.310 1.160 ;
        RECT  13.970 0.820 14.200 4.180 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.260 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.250 -0.400 13.590 1.005 ;
        RECT  11.275 -0.400 11.615 0.880 ;
        RECT  6.295 -0.400 6.635 0.950 ;
        RECT  1.210 -0.400 1.550 1.450 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.250 3.330 13.590 5.280 ;
        RECT  11.990 4.200 12.330 5.280 ;
        RECT  10.415 3.665 10.755 5.280 ;
        RECT  7.815 3.480 8.155 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.215 ;
        RECT  0.170 1.985 2.445 2.215 ;
        RECT  2.160 1.985 2.445 2.325 ;
        RECT  0.170 0.645 0.400 3.360 ;
        RECT  0.170 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 0.970 2.785 ;
        RECT  0.630 2.520 1.985 2.785 ;
        RECT  1.755 2.520 1.985 3.340 ;
        RECT  1.755 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  1.970 0.630 5.105 0.860 ;
        RECT  4.795 0.630 5.105 1.375 ;
        RECT  1.970 0.630 2.310 1.450 ;
        RECT  7.325 1.240 7.665 1.580 ;
        RECT  7.380 1.240 7.665 2.690 ;
        RECT  7.380 2.460 8.830 2.690 ;
        RECT  8.490 2.460 8.830 2.800 ;
        RECT  3.520 2.285 3.845 3.115 ;
        RECT  7.275 2.720 7.615 3.295 ;
        RECT  3.520 2.885 5.105 3.115 ;
        RECT  7.380 1.240 7.615 3.295 ;
        RECT  4.875 3.065 7.615 3.295 ;
        RECT  6.865 0.780 8.125 1.010 ;
        RECT  5.335 1.070 5.875 1.410 ;
        RECT  5.335 1.180 7.095 1.410 ;
        RECT  6.865 0.780 7.095 2.100 ;
        RECT  6.780 1.180 7.095 2.100 ;
        RECT  3.135 1.555 4.305 1.785 ;
        RECT  7.895 0.780 8.125 2.020 ;
        RECT  3.135 1.555 3.420 1.895 ;
        RECT  7.895 1.790 9.290 2.020 ;
        RECT  6.780 1.760 7.120 2.100 ;
        RECT  8.615 1.790 9.290 2.130 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  4.075 2.290 4.530 2.655 ;
        RECT  5.335 1.070 5.565 2.835 ;
        RECT  4.075 2.425 5.565 2.655 ;
        RECT  5.335 2.550 6.040 2.835 ;
        RECT  9.060 1.790 9.290 3.240 ;
        RECT  9.060 2.900 9.590 3.240 ;
        RECT  8.355 0.630 10.810 0.860 ;
        RECT  10.470 0.630 10.810 0.950 ;
        RECT  8.355 0.630 8.695 0.970 ;
        RECT  9.135 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  9.625 1.970 10.150 2.200 ;
        RECT  11.470 2.650 12.050 2.940 ;
        RECT  9.920 2.860 11.700 3.200 ;
        RECT  9.920 1.970 10.150 3.710 ;
        RECT  8.970 3.480 10.150 3.710 ;
        RECT  8.970 3.480 9.310 3.820 ;
        RECT  10.085 1.180 12.340 1.410 ;
        RECT  10.085 1.180 10.425 1.720 ;
        RECT  12.110 1.180 12.340 1.925 ;
        RECT  12.330 1.695 12.830 2.555 ;
        RECT  12.330 2.160 12.985 2.555 ;
        RECT  12.330 1.695 12.560 3.400 ;
        RECT  12.030 3.170 12.560 3.400 ;
        RECT  12.030 3.170 12.260 3.895 ;
        RECT  11.190 3.665 12.260 3.895 ;
        RECT  11.190 3.665 11.530 4.005 ;
        RECT  0.170 1.985 1.60 2.215 ;
        RECT  1.970 0.630 4.60 0.860 ;
        RECT  4.875 3.065 6.30 3.295 ;
        RECT  8.355 0.630 9.20 0.860 ;
        RECT  10.085 1.180 11.40 1.410 ;
    END
END DFFRSX1

MACRO DFFRSX0
    CLASS CORE ;
    FOREIGN DFFRSX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.592  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.065 2.860 12.625 3.350 ;
        RECT  12.395 0.630 12.625 3.350 ;
        RECT  11.730 0.630 12.625 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.380 2.235 4.915 2.695 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.250 10.220 2.760 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.248  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.660 2.250 11.215 2.845 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.443  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.965 2.860 13.735 3.240 ;
        RECT  12.855 3.010 13.195 3.350 ;
        RECT  12.965 1.170 13.195 3.350 ;
        RECT  12.855 1.170 13.195 1.510 ;
        END
    END QN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.605 2.160 6.175 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.120 3.810 13.040 5.280 ;
        RECT  9.565 3.910 9.900 5.280 ;
        RECT  6.970 3.630 7.310 5.280 ;
        RECT  4.810 3.910 6.085 5.280 ;
        RECT  1.470 3.520 2.335 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.865 -0.400 13.205 0.710 ;
        RECT  10.700 -0.400 11.040 0.950 ;
        RECT  6.030 -0.400 6.315 1.400 ;
        RECT  1.100 -0.400 1.440 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.970 ;
        RECT  0.115 1.740 2.335 1.970 ;
        RECT  2.050 1.740 2.335 2.460 ;
        RECT  0.115 0.630 0.345 3.060 ;
        RECT  0.115 2.770 1.010 3.060 ;
        RECT  2.565 1.285 3.470 1.545 ;
        RECT  0.575 2.200 1.565 2.540 ;
        RECT  1.335 2.200 1.565 3.060 ;
        RECT  1.335 2.690 2.795 3.060 ;
        RECT  2.565 1.285 2.795 4.140 ;
        RECT  2.565 3.910 3.810 4.140 ;
        RECT  3.470 3.910 3.810 4.250 ;
        RECT  1.900 0.825 4.870 1.055 ;
        RECT  1.900 0.825 2.240 1.510 ;
        RECT  4.530 0.825 4.870 1.545 ;
        RECT  7.005 1.230 7.265 1.570 ;
        RECT  7.035 1.230 7.265 3.200 ;
        RECT  3.190 2.840 3.530 3.180 ;
        RECT  6.510 2.860 8.260 3.200 ;
        RECT  3.300 2.840 3.530 3.675 ;
        RECT  6.510 2.860 6.740 3.675 ;
        RECT  3.300 3.445 6.740 3.675 ;
        RECT  6.545 0.765 7.725 0.995 ;
        RECT  5.145 1.230 5.570 1.905 ;
        RECT  5.145 1.675 6.775 1.905 ;
        RECT  3.025 1.775 5.375 2.005 ;
        RECT  6.545 0.765 6.775 2.110 ;
        RECT  6.405 1.675 6.775 2.110 ;
        RECT  3.025 1.775 4.090 2.180 ;
        RECT  7.495 0.765 7.725 2.485 ;
        RECT  7.495 2.190 8.875 2.485 ;
        RECT  3.860 1.775 4.090 3.180 ;
        RECT  5.145 1.230 5.375 3.200 ;
        RECT  3.860 2.840 4.200 3.180 ;
        RECT  5.145 2.860 5.485 3.200 ;
        RECT  8.590 2.190 8.875 3.435 ;
        RECT  7.955 0.630 10.170 0.860 ;
        RECT  7.955 0.630 8.240 0.970 ;
        RECT  9.830 0.630 10.170 0.970 ;
        RECT  8.800 1.170 9.140 1.510 ;
        RECT  10.140 3.075 10.500 3.525 ;
        RECT  10.140 3.125 11.375 3.525 ;
        RECT  9.105 3.285 11.375 3.525 ;
        RECT  9.105 1.280 9.335 3.970 ;
        RECT  8.270 3.665 9.335 3.970 ;
        RECT  11.730 1.310 12.070 2.170 ;
        RECT  9.750 1.690 12.070 1.920 ;
        RECT  9.750 1.690 10.090 2.020 ;
        RECT  11.605 1.830 12.165 2.170 ;
        RECT  11.605 1.690 11.835 4.155 ;
        RECT  10.695 3.925 11.835 4.155 ;
        RECT  10.695 3.925 11.035 4.250 ;
        RECT  0.115 1.740 1.80 1.970 ;
        RECT  1.900 0.825 3.40 1.055 ;
        RECT  3.300 3.445 5.90 3.675 ;
        RECT  3.025 1.775 4.50 2.005 ;
        RECT  7.955 0.630 9.60 0.860 ;
        RECT  9.105 3.285 10.80 3.525 ;
        RECT  9.750 1.690 11.50 1.920 ;
    END
END DFFRSX0

MACRO DFFRSQX4
    CLASS CORE ;
    FOREIGN DFFRSQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.198  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  17.120 1.240 17.460 4.030 ;
        RECT  15.800 2.250 17.460 2.630 ;
        RECT  15.800 0.790 16.140 2.630 ;
        RECT  15.680 2.790 16.030 4.030 ;
        RECT  15.800 0.790 16.030 4.030 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.511  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.905 1.640 14.365 2.560 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.655 2.230 13.265 2.630 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.600 1.660 8.065 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.640 0.400 ;
        RECT  16.560 -0.400 16.900 0.720 ;
        RECT  15.040 -0.400 15.380 0.835 ;
        RECT  13.430 -0.400 13.770 0.710 ;
        RECT  7.830 -0.400 8.115 0.970 ;
        RECT  2.255 -0.400 3.825 0.665 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.640 5.280 ;
        RECT  16.400 2.860 16.740 5.280 ;
        RECT  14.875 4.060 15.215 5.280 ;
        RECT  12.435 3.910 13.895 5.280 ;
        RECT  10.135 3.965 10.475 5.280 ;
        RECT  7.715 2.910 8.015 5.280 ;
        RECT  2.410 3.965 3.845 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.765 1.815 2.105 2.095 ;
        RECT  1.375 1.860 4.020 2.095 ;
        RECT  3.790 1.860 4.020 2.800 ;
        RECT  3.790 2.460 4.130 2.800 ;
        RECT  1.375 1.860 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.965 1.355 4.535 1.585 ;
        RECT  0.965 1.290 1.305 1.630 ;
        RECT  2.925 1.355 4.535 1.630 ;
        RECT  4.245 1.355 4.535 1.695 ;
        RECT  5.475 1.160 5.810 1.500 ;
        RECT  4.765 1.270 5.810 1.500 ;
        RECT  1.835 2.325 3.180 2.665 ;
        RECT  2.840 2.325 3.180 3.275 ;
        RECT  4.765 1.270 4.995 3.540 ;
        RECT  2.840 3.045 4.995 3.275 ;
        RECT  4.735 3.200 5.080 3.540 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.505 4.415 3.735 ;
        RECT  4.185 3.505 4.415 4.000 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  5.500 2.980 5.840 4.000 ;
        RECT  4.185 3.770 5.840 4.000 ;
        RECT  0.365 0.640 0.705 1.015 ;
        RECT  4.120 0.630 6.270 0.860 ;
        RECT  0.365 0.785 2.025 1.015 ;
        RECT  4.120 0.630 4.350 1.125 ;
        RECT  1.795 0.895 4.350 1.125 ;
        RECT  6.040 0.630 6.270 1.605 ;
        RECT  6.040 1.320 6.625 1.605 ;
        RECT  8.345 0.775 9.495 1.005 ;
        RECT  6.500 0.735 7.370 1.090 ;
        RECT  7.140 1.200 8.575 1.430 ;
        RECT  9.265 0.775 9.495 2.090 ;
        RECT  9.265 1.860 10.930 2.090 ;
        RECT  8.345 0.775 8.575 2.100 ;
        RECT  8.295 1.200 8.575 2.100 ;
        RECT  7.140 0.735 7.370 2.150 ;
        RECT  6.795 1.920 7.370 2.150 ;
        RECT  10.590 1.860 10.930 2.200 ;
        RECT  6.795 1.920 7.025 3.195 ;
        RECT  6.685 2.855 7.025 3.195 ;
        RECT  11.260 1.670 11.600 2.010 ;
        RECT  5.225 1.835 6.455 2.120 ;
        RECT  8.805 1.240 9.035 2.680 ;
        RECT  8.805 2.340 9.505 2.680 ;
        RECT  11.260 1.670 11.490 2.680 ;
        RECT  7.255 2.450 11.490 2.680 ;
        RECT  8.395 2.450 8.735 2.860 ;
        RECT  6.225 1.835 6.455 3.655 ;
        RECT  8.395 2.450 8.625 3.855 ;
        RECT  7.255 2.450 7.485 3.655 ;
        RECT  6.225 3.425 7.485 3.655 ;
        RECT  9.605 3.505 11.115 3.735 ;
        RECT  10.885 3.505 11.115 4.100 ;
        RECT  8.395 3.625 9.835 3.855 ;
        RECT  10.885 3.760 11.225 4.100 ;
        RECT  9.725 0.630 12.965 0.860 ;
        RECT  12.155 0.630 12.965 0.950 ;
        RECT  9.725 0.630 10.020 1.500 ;
        RECT  10.830 1.100 11.170 1.440 ;
        RECT  10.830 1.210 12.060 1.440 ;
        RECT  11.830 1.210 12.060 3.275 ;
        RECT  12.995 2.860 14.890 3.090 ;
        RECT  14.595 2.270 14.890 3.090 ;
        RECT  8.945 3.045 13.335 3.275 ;
        RECT  8.945 3.045 9.285 3.395 ;
        RECT  11.455 3.045 11.745 3.980 ;
        RECT  14.415 1.110 14.825 1.410 ;
        RECT  12.290 1.180 14.825 1.410 ;
        RECT  14.435 1.110 14.825 1.420 ;
        RECT  12.290 1.180 12.630 1.675 ;
        RECT  14.595 1.110 14.825 2.040 ;
        RECT  14.595 1.810 15.350 2.040 ;
        RECT  15.120 1.810 15.350 3.550 ;
        RECT  14.315 3.320 15.350 3.550 ;
        RECT  14.315 3.320 14.655 3.660 ;
        RECT  1.375 1.860 3.70 2.095 ;
        RECT  0.965 1.355 3.70 1.585 ;
        RECT  2.840 3.045 3.30 3.275 ;
        RECT  2.030 3.505 3.20 3.735 ;
        RECT  0.180 3.600 1.60 3.830 ;
        RECT  4.120 0.630 5.80 0.860 ;
        RECT  1.795 0.895 3.90 1.125 ;
        RECT  7.255 2.450 10.50 2.680 ;
        RECT  9.725 0.630 11.60 0.860 ;
        RECT  8.945 3.045 12.70 3.275 ;
        RECT  12.290 1.180 13.60 1.410 ;
    END
END DFFRSQX4

MACRO DFFRSQX2
    CLASS CORE ;
    FOREIGN DFFRSQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.355 1.240 13.750 3.550 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.780 2.070 11.225 2.630 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.358  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.640 11.845 2.585 ;
        END
    END SN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.820 1.640 5.105 2.100 ;
        RECT  4.535 1.640 5.105 2.020 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.290 2.140 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  12.850 3.950 14.310 5.280 ;
        RECT  11.370 3.730 11.710 5.280 ;
        RECT  10.000 3.910 10.340 5.280 ;
        RECT  7.730 3.480 8.070 5.280 ;
        RECT  6.430 3.525 6.770 5.280 ;
        RECT  5.130 3.525 5.470 5.280 ;
        RECT  1.500 3.805 2.900 5.280 ;
        RECT  0.180 3.780 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  12.850 -0.400 14.310 0.720 ;
        RECT  11.155 -0.400 11.495 0.950 ;
        RECT  6.060 -0.400 6.400 0.950 ;
        RECT  1.210 -0.400 1.550 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.360 0.520 2.070 ;
        RECT  0.130 1.840 2.405 2.070 ;
        RECT  2.120 1.840 2.405 2.490 ;
        RECT  0.130 1.360 0.360 3.100 ;
        RECT  0.130 2.870 1.080 3.100 ;
        RECT  0.740 2.870 1.080 3.160 ;
        RECT  2.635 1.090 3.540 1.325 ;
        RECT  0.590 2.300 0.930 2.640 ;
        RECT  0.590 2.410 1.630 2.640 ;
        RECT  1.400 2.410 1.630 3.190 ;
        RECT  1.400 2.850 2.865 3.190 ;
        RECT  2.635 1.090 2.865 3.575 ;
        RECT  2.635 3.345 3.930 3.575 ;
        RECT  3.590 3.345 3.930 3.820 ;
        RECT  1.970 0.630 4.940 0.860 ;
        RECT  4.600 0.630 4.940 1.370 ;
        RECT  1.970 0.630 2.310 1.530 ;
        RECT  7.090 1.240 7.380 1.580 ;
        RECT  7.150 1.240 7.380 3.295 ;
        RECT  7.150 2.320 8.865 2.550 ;
        RECT  8.525 2.320 8.865 2.660 ;
        RECT  3.510 2.310 3.845 3.115 ;
        RECT  3.510 2.885 5.105 3.115 ;
        RECT  7.150 2.320 7.530 3.295 ;
        RECT  4.875 3.065 7.530 3.295 ;
        RECT  6.630 0.780 7.840 1.010 ;
        RECT  5.300 1.070 5.640 1.410 ;
        RECT  5.300 1.180 6.860 1.410 ;
        RECT  3.095 1.555 3.390 1.895 ;
        RECT  7.610 0.780 7.840 1.940 ;
        RECT  6.630 0.780 6.860 2.175 ;
        RECT  3.095 1.665 4.305 1.895 ;
        RECT  7.610 1.710 8.385 1.940 ;
        RECT  8.045 1.820 9.325 2.050 ;
        RECT  6.580 1.840 6.920 2.175 ;
        RECT  4.075 1.665 4.305 2.655 ;
        RECT  4.075 2.290 4.520 2.655 ;
        RECT  5.335 1.070 5.565 2.835 ;
        RECT  4.075 2.425 5.565 2.655 ;
        RECT  9.095 1.820 9.325 3.080 ;
        RECT  5.335 2.550 6.010 2.835 ;
        RECT  9.095 2.740 9.590 3.080 ;
        RECT  8.070 0.630 10.735 0.860 ;
        RECT  8.070 0.630 8.355 0.970 ;
        RECT  10.395 0.630 10.735 1.040 ;
        RECT  9.165 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  12.320 2.750 12.660 3.090 ;
        RECT  9.820 2.860 12.660 3.090 ;
        RECT  10.760 2.860 11.100 3.200 ;
        RECT  9.820 1.970 10.050 3.550 ;
        RECT  8.950 3.320 10.050 3.550 ;
        RECT  8.950 3.320 9.290 3.660 ;
        RECT  11.985 0.630 12.325 1.410 ;
        RECT  10.985 1.180 13.120 1.410 ;
        RECT  10.115 1.400 11.215 1.630 ;
        RECT  10.115 1.400 10.455 1.740 ;
        RECT  12.890 1.180 13.120 3.720 ;
        RECT  12.090 3.490 13.120 3.720 ;
        RECT  12.090 3.490 12.430 4.060 ;
        RECT  0.130 1.840 1.90 2.070 ;
        RECT  1.970 0.630 3.70 0.860 ;
        RECT  4.875 3.065 6.60 3.295 ;
        RECT  8.070 0.630 9.70 0.860 ;
        RECT  9.820 2.860 11.60 3.090 ;
        RECT  10.985 1.180 12.80 1.410 ;
    END
END DFFRSQX2

MACRO DFFRSQX1
    CLASS CORE ;
    FOREIGN DFFRSQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.105 2.025 ;
        END
    END D
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.270  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.465 1.640 11.845 2.305 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.835 2.045 11.215 2.630 ;
        RECT  10.520 2.045 11.215 2.385 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.712  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.880 2.400 13.735 2.630 ;
        RECT  13.355 2.250 13.735 2.630 ;
        RECT  13.355 1.235 13.585 2.630 ;
        RECT  12.730 1.235 13.585 1.465 ;
        RECT  12.620 3.635 13.110 3.920 ;
        RECT  12.880 2.400 13.110 3.920 ;
        RECT  12.730 0.700 12.960 1.465 ;
        RECT  12.655 3.615 13.110 3.920 ;
        RECT  12.620 0.700 12.960 1.040 ;
        END
    END Q
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.335 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  13.340 -0.400 13.680 1.005 ;
        RECT  11.275 -0.400 11.615 0.880 ;
        RECT  6.295 -0.400 6.635 0.925 ;
        RECT  1.210 -0.400 1.550 1.450 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  13.340 3.330 13.680 5.280 ;
        RECT  11.990 4.170 12.330 5.280 ;
        RECT  10.415 3.665 10.755 5.280 ;
        RECT  7.815 3.480 8.155 5.280 ;
        RECT  6.515 3.525 6.855 5.280 ;
        RECT  5.200 3.525 5.540 5.280 ;
        RECT  1.540 3.840 2.820 5.280 ;
        RECT  0.180 3.840 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.645 0.520 2.215 ;
        RECT  0.170 1.985 2.445 2.215 ;
        RECT  2.160 1.985 2.445 2.325 ;
        RECT  0.170 0.645 0.400 3.360 ;
        RECT  0.170 3.020 1.120 3.360 ;
        RECT  2.675 1.090 3.570 1.325 ;
        RECT  0.630 2.445 0.970 2.785 ;
        RECT  0.630 2.520 1.985 2.785 ;
        RECT  1.755 2.520 1.985 3.340 ;
        RECT  1.755 3.000 2.905 3.340 ;
        RECT  2.675 1.090 2.905 3.575 ;
        RECT  2.675 3.345 4.140 3.575 ;
        RECT  3.800 3.345 4.140 3.665 ;
        RECT  1.970 0.630 5.105 0.860 ;
        RECT  4.795 0.630 5.105 1.410 ;
        RECT  1.970 0.630 2.310 1.450 ;
        RECT  7.325 1.240 7.665 1.580 ;
        RECT  7.380 1.240 7.665 2.690 ;
        RECT  7.380 2.460 8.830 2.690 ;
        RECT  8.490 2.460 8.830 2.800 ;
        RECT  3.520 2.295 3.845 3.115 ;
        RECT  7.265 2.720 7.615 3.295 ;
        RECT  3.520 2.885 5.105 3.115 ;
        RECT  7.380 1.240 7.615 3.295 ;
        RECT  4.875 3.065 7.615 3.295 ;
        RECT  6.865 0.780 8.125 1.010 ;
        RECT  5.335 1.070 5.875 1.385 ;
        RECT  6.865 0.780 7.095 1.385 ;
        RECT  5.335 1.155 7.095 1.385 ;
        RECT  5.335 1.070 5.870 1.410 ;
        RECT  3.135 1.555 4.305 1.785 ;
        RECT  7.895 0.780 8.125 2.020 ;
        RECT  3.135 1.555 3.420 1.895 ;
        RECT  6.780 1.155 7.010 2.360 ;
        RECT  7.895 1.790 9.290 2.020 ;
        RECT  8.775 1.790 9.290 2.130 ;
        RECT  4.075 1.555 4.305 2.655 ;
        RECT  6.780 2.020 7.120 2.360 ;
        RECT  4.075 2.290 4.530 2.655 ;
        RECT  5.335 1.070 5.565 2.835 ;
        RECT  4.075 2.425 5.565 2.655 ;
        RECT  5.335 2.550 6.040 2.835 ;
        RECT  9.060 1.790 9.290 3.130 ;
        RECT  9.250 2.900 9.590 3.240 ;
        RECT  8.355 0.630 10.810 0.860 ;
        RECT  10.470 0.630 10.810 0.950 ;
        RECT  8.355 0.630 8.695 0.970 ;
        RECT  9.135 1.170 9.855 1.510 ;
        RECT  9.625 1.170 9.855 2.200 ;
        RECT  9.625 1.970 10.150 2.200 ;
        RECT  11.470 2.635 12.050 2.945 ;
        RECT  9.920 2.860 11.700 3.200 ;
        RECT  9.920 1.970 10.150 3.710 ;
        RECT  8.970 3.480 10.150 3.710 ;
        RECT  8.970 3.480 9.310 3.820 ;
        RECT  10.085 1.180 12.340 1.410 ;
        RECT  10.085 1.180 10.425 1.730 ;
        RECT  12.110 1.180 12.340 1.925 ;
        RECT  12.330 1.695 12.940 1.980 ;
        RECT  12.330 1.695 12.560 3.405 ;
        RECT  12.030 3.175 12.560 3.405 ;
        RECT  12.030 3.175 12.260 3.895 ;
        RECT  11.190 3.665 12.260 3.895 ;
        RECT  11.190 3.665 11.530 4.005 ;
        RECT  0.170 1.985 1.30 2.215 ;
        RECT  1.970 0.630 4.40 0.860 ;
        RECT  4.875 3.065 6.60 3.295 ;
        RECT  8.355 0.630 9.70 0.860 ;
        RECT  10.085 1.180 11.60 1.410 ;
    END
END DFFRSQX1

MACRO DFFRSQX0
    CLASS CORE ;
    FOREIGN DFFRSQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.592  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.065 2.860 12.485 3.350 ;
        RECT  12.255 0.630 12.485 3.350 ;
        RECT  11.730 0.630 12.485 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.380 2.235 4.915 2.695 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.575 2.250 10.220 2.760 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.248  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.660 2.250 11.215 2.845 ;
        END
    END SN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.605 2.135 6.175 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  12.080 3.810 12.420 5.280 ;
        RECT  9.565 3.910 9.900 5.280 ;
        RECT  6.970 3.630 7.310 5.280 ;
        RECT  4.810 3.910 6.085 5.280 ;
        RECT  1.470 3.520 2.335 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  10.700 -0.400 11.040 0.950 ;
        RECT  6.030 -0.400 6.315 1.400 ;
        RECT  1.100 -0.400 1.440 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.630 0.520 1.970 ;
        RECT  0.115 1.740 2.335 1.970 ;
        RECT  2.050 1.740 2.335 2.460 ;
        RECT  0.115 0.630 0.345 3.060 ;
        RECT  0.115 2.770 1.010 3.060 ;
        RECT  2.565 1.285 3.470 1.545 ;
        RECT  0.575 2.200 1.565 2.540 ;
        RECT  1.335 2.200 1.565 3.060 ;
        RECT  1.335 2.690 2.795 3.060 ;
        RECT  2.565 1.285 2.795 4.140 ;
        RECT  2.565 3.910 3.810 4.140 ;
        RECT  3.470 3.910 3.810 4.250 ;
        RECT  1.900 0.825 4.870 1.055 ;
        RECT  1.900 0.825 2.240 1.510 ;
        RECT  4.530 0.825 4.870 1.545 ;
        RECT  7.005 1.230 7.265 1.570 ;
        RECT  7.035 1.230 7.265 3.200 ;
        RECT  3.190 2.840 3.530 3.180 ;
        RECT  6.510 2.860 8.260 3.200 ;
        RECT  3.300 2.840 3.530 3.675 ;
        RECT  6.510 2.860 6.740 3.675 ;
        RECT  3.300 3.445 6.740 3.675 ;
        RECT  6.545 0.765 7.725 0.995 ;
        RECT  5.145 1.230 5.570 1.905 ;
        RECT  5.145 1.675 6.775 1.905 ;
        RECT  3.025 1.775 5.375 2.005 ;
        RECT  6.545 0.765 6.775 2.110 ;
        RECT  6.405 1.675 6.775 2.110 ;
        RECT  3.025 1.775 4.090 2.180 ;
        RECT  7.495 0.765 7.725 2.485 ;
        RECT  7.495 2.190 8.875 2.485 ;
        RECT  3.860 1.775 4.090 3.180 ;
        RECT  5.145 1.230 5.375 3.200 ;
        RECT  3.860 2.840 4.200 3.180 ;
        RECT  5.145 2.860 5.485 3.200 ;
        RECT  8.590 2.190 8.875 3.435 ;
        RECT  7.955 0.630 10.170 0.860 ;
        RECT  7.955 0.630 8.240 0.970 ;
        RECT  9.830 0.630 10.170 0.970 ;
        RECT  8.800 1.170 9.140 1.510 ;
        RECT  10.140 3.075 10.500 3.525 ;
        RECT  9.105 3.125 11.375 3.525 ;
        RECT  9.105 1.280 9.335 3.970 ;
        RECT  8.270 3.665 9.335 3.970 ;
        RECT  9.750 1.310 12.025 1.540 ;
        RECT  11.605 1.310 12.025 1.650 ;
        RECT  9.750 1.310 10.090 2.020 ;
        RECT  11.605 1.310 11.835 4.155 ;
        RECT  10.695 3.925 11.835 4.155 ;
        RECT  10.695 3.925 11.035 4.250 ;
        RECT  0.115 1.740 1.60 1.970 ;
        RECT  1.900 0.825 3.90 1.055 ;
        RECT  3.300 3.445 5.70 3.675 ;
        RECT  3.025 1.775 4.00 2.005 ;
        RECT  7.955 0.630 9.30 0.860 ;
        RECT  9.105 3.125 10.20 3.525 ;
        RECT  9.750 1.310 11.70 1.540 ;
    END
END DFFRSQX0

MACRO DFFRQX4
    CLASS CORE ;
    FOREIGN DFFRQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 2.075 16.885 3.880 ;
        RECT  14.330 2.075 16.885 2.305 ;
        RECT  15.770 1.130 16.110 2.305 ;
        RECT  15.050 2.075 15.390 3.880 ;
        RECT  14.330 1.130 14.670 2.305 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.844  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.290 1.640 13.105 2.020 ;
        RECT  12.290 1.640 12.630 2.190 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.760 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.715 1.660 7.435 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 1.470 ;
        RECT  15.050 -0.400 15.390 1.470 ;
        RECT  12.800 -0.400 13.140 0.950 ;
        RECT  7.230 -0.400 7.515 0.970 ;
        RECT  1.750 -0.400 3.225 0.655 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 2.640 16.110 5.280 ;
        RECT  14.330 2.640 14.670 5.280 ;
        RECT  11.490 3.760 12.950 5.280 ;
        RECT  9.315 4.170 9.655 5.280 ;
        RECT  6.825 3.925 7.165 5.280 ;
        RECT  2.410 3.985 3.245 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.805 1.920 2.090 ;
        RECT  1.375 1.860 3.420 2.090 ;
        RECT  3.190 1.860 3.420 2.800 ;
        RECT  3.190 2.460 3.530 2.800 ;
        RECT  1.375 1.805 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  0.780 1.345 3.935 1.575 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  2.325 1.345 3.935 1.630 ;
        RECT  3.645 1.345 3.935 1.695 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  2.030 3.525 5.200 3.755 ;
        RECT  4.860 3.010 5.200 3.755 ;
        RECT  0.180 3.600 2.220 3.830 ;
        RECT  4.875 1.160 5.210 1.500 ;
        RECT  4.165 1.270 5.210 1.500 ;
        RECT  1.835 2.325 2.580 2.665 ;
        RECT  4.165 1.270 4.395 3.295 ;
        RECT  2.240 2.325 2.580 3.295 ;
        RECT  4.140 2.955 4.480 3.295 ;
        RECT  2.240 3.065 4.480 3.295 ;
        RECT  0.180 0.640 0.520 1.015 ;
        RECT  3.520 0.700 5.670 0.930 ;
        RECT  0.180 0.785 1.520 1.015 ;
        RECT  1.290 0.885 3.750 1.115 ;
        RECT  5.440 0.700 5.670 1.660 ;
        RECT  5.440 1.320 6.025 1.660 ;
        RECT  7.745 0.775 8.895 1.005 ;
        RECT  5.900 0.735 6.770 1.090 ;
        RECT  6.255 0.735 6.770 1.430 ;
        RECT  6.255 1.200 7.975 1.430 ;
        RECT  8.665 0.775 8.895 2.090 ;
        RECT  8.665 1.860 10.330 2.090 ;
        RECT  6.255 0.735 6.485 2.150 ;
        RECT  9.990 1.860 10.330 2.200 ;
        RECT  7.745 0.775 7.975 2.225 ;
        RECT  7.665 1.200 7.975 2.225 ;
        RECT  6.050 1.920 6.390 3.235 ;
        RECT  4.625 1.820 4.935 2.120 ;
        RECT  10.660 1.670 10.945 2.010 ;
        RECT  4.625 1.890 5.810 2.120 ;
        RECT  8.205 1.240 8.435 2.805 ;
        RECT  8.205 2.340 8.685 2.805 ;
        RECT  8.205 2.520 10.890 2.805 ;
        RECT  10.660 1.670 10.890 2.805 ;
        RECT  7.585 2.575 10.890 2.805 ;
        RECT  7.585 2.575 7.925 2.915 ;
        RECT  5.470 1.890 5.810 3.695 ;
        RECT  5.470 3.465 7.815 3.695 ;
        RECT  7.585 2.575 7.815 3.940 ;
        RECT  7.585 3.710 10.170 3.940 ;
        RECT  9.940 3.710 10.170 4.250 ;
        RECT  9.940 3.965 10.280 4.250 ;
        RECT  9.125 0.630 12.340 0.860 ;
        RECT  11.530 0.630 12.340 0.950 ;
        RECT  9.125 0.630 9.420 1.500 ;
        RECT  10.230 1.100 10.570 1.440 ;
        RECT  10.230 1.210 11.405 1.440 ;
        RECT  11.175 1.210 11.405 3.395 ;
        RECT  13.295 2.150 13.600 2.650 ;
        RECT  13.315 2.120 13.600 2.650 ;
        RECT  11.175 2.420 13.600 2.650 ;
        RECT  12.050 2.420 12.390 3.150 ;
        RECT  11.175 2.420 11.460 3.395 ;
        RECT  8.125 3.165 11.460 3.395 ;
        RECT  8.125 3.165 8.465 3.480 ;
        RECT  10.485 3.165 10.800 3.860 ;
        RECT  10.510 3.165 10.800 3.890 ;
        RECT  11.635 1.180 14.060 1.410 ;
        RECT  13.560 1.180 14.060 1.520 ;
        RECT  11.635 1.180 11.975 1.675 ;
        RECT  13.830 1.180 14.060 3.240 ;
        RECT  13.570 3.010 13.910 3.880 ;
        RECT  1.375 1.860 2.70 2.090 ;
        RECT  0.780 1.345 2.60 1.575 ;
        RECT  2.030 3.525 4.50 3.755 ;
        RECT  0.180 3.600 1.80 3.830 ;
        RECT  2.240 3.065 3.20 3.295 ;
        RECT  3.520 0.700 4.30 0.930 ;
        RECT  1.290 0.885 2.20 1.115 ;
        RECT  8.205 2.520 9.50 2.805 ;
        RECT  7.585 2.575 9.10 2.805 ;
        RECT  5.470 3.465 6.40 3.695 ;
        RECT  7.585 3.710 9.80 3.940 ;
        RECT  9.125 0.630 11.40 0.860 ;
        RECT  11.175 2.420 12.40 2.650 ;
        RECT  8.125 3.165 10.30 3.395 ;
        RECT  11.635 1.180 13.20 1.410 ;
    END
END DFFRQX4

MACRO DFFRQX2
    CLASS CORE ;
    FOREIGN DFFRQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.230 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.095 1.240 12.490 3.550 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.524  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.045 2.220 10.605 2.680 ;
        END
    END RN
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.400 1.640 4.915 2.120 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.650 5.560 2.195 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.230 5.280 ;
        RECT  11.590 3.950 13.050 5.280 ;
        RECT  9.620 4.170 9.960 5.280 ;
        RECT  7.200 3.660 7.540 5.280 ;
        RECT  5.900 3.525 6.240 5.280 ;
        RECT  4.600 3.525 4.940 5.280 ;
        RECT  1.470 3.805 2.400 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.230 0.400 ;
        RECT  11.590 -0.400 13.050 0.720 ;
        RECT  10.230 -0.400 10.570 1.040 ;
        RECT  5.390 -0.400 5.730 0.925 ;
        RECT  0.780 -0.400 1.120 1.050 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.360 0.520 2.510 ;
        RECT  0.115 2.280 1.905 2.510 ;
        RECT  1.620 2.280 1.905 2.620 ;
        RECT  0.115 2.280 0.345 4.070 ;
        RECT  0.115 3.730 0.620 4.070 ;
        RECT  2.135 1.305 3.040 1.645 ;
        RECT  0.575 2.850 2.365 3.190 ;
        RECT  2.135 1.305 2.365 3.575 ;
        RECT  2.135 3.345 3.630 3.575 ;
        RECT  3.290 3.345 3.630 3.685 ;
        RECT  1.580 0.630 4.240 0.950 ;
        RECT  1.580 0.630 1.920 1.090 ;
        RECT  6.420 1.240 6.710 1.845 ;
        RECT  6.620 1.615 6.850 3.295 ;
        RECT  7.920 2.360 8.260 2.700 ;
        RECT  6.620 2.470 8.260 2.700 ;
        RECT  3.010 2.505 3.350 3.115 ;
        RECT  3.010 2.885 4.910 3.115 ;
        RECT  6.620 2.470 7.000 3.295 ;
        RECT  4.680 3.065 7.000 3.295 ;
        RECT  5.960 0.780 7.310 1.010 ;
        RECT  4.630 1.155 6.190 1.385 ;
        RECT  5.960 0.780 6.190 1.385 ;
        RECT  4.630 1.070 4.970 1.410 ;
        RECT  3.680 1.180 4.970 1.410 ;
        RECT  7.080 0.780 7.310 1.980 ;
        RECT  7.080 1.750 7.660 1.980 ;
        RECT  7.320 1.900 8.740 2.130 ;
        RECT  2.595 1.880 3.910 2.220 ;
        RECT  3.680 1.180 3.910 2.655 ;
        RECT  6.050 2.075 6.390 2.375 ;
        RECT  3.680 2.315 4.020 2.655 ;
        RECT  6.050 2.075 6.280 2.655 ;
        RECT  3.680 2.425 6.280 2.655 ;
        RECT  8.510 1.900 8.740 3.130 ;
        RECT  5.140 2.425 5.480 2.835 ;
        RECT  8.510 2.790 9.010 3.130 ;
        RECT  7.540 0.630 9.810 0.970 ;
        RECT  9.470 0.630 9.810 1.040 ;
        RECT  8.440 1.330 9.200 1.670 ;
        RECT  8.970 1.330 9.200 2.560 ;
        RECT  8.970 2.330 9.470 2.560 ;
        RECT  9.240 2.915 11.135 3.145 ;
        RECT  10.180 2.915 11.135 3.260 ;
        RECT  10.180 2.915 10.520 3.440 ;
        RECT  9.240 2.330 9.470 3.715 ;
        RECT  8.385 3.485 9.470 3.715 ;
        RECT  8.385 3.485 8.725 3.825 ;
        RECT  10.795 1.360 11.135 1.990 ;
        RECT  9.430 1.760 11.595 1.990 ;
        RECT  9.430 1.760 9.730 2.100 ;
        RECT  11.365 1.760 11.595 3.720 ;
        RECT  10.940 3.490 11.595 3.720 ;
        RECT  10.940 3.490 11.170 4.180 ;
        RECT  10.830 3.840 11.170 4.180 ;
        RECT  1.580 0.630 3.50 0.950 ;
        RECT  4.680 3.065 6.00 3.295 ;
        RECT  3.680 2.425 5.40 2.655 ;
        RECT  7.540 0.630 8.80 0.970 ;
        RECT  9.430 1.760 10.40 1.990 ;
    END
END DFFRQX2

MACRO DFFRQX1
    CLASS CORE ;
    FOREIGN DFFRQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.655 2.025 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.403  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.050 1.640 10.610 2.085 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.680  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.620 2.400 12.475 2.630 ;
        RECT  11.860 2.250 12.475 2.630 ;
        RECT  11.860 1.235 12.090 2.630 ;
        RECT  11.360 1.235 12.090 1.465 ;
        RECT  11.360 3.435 11.850 3.720 ;
        RECT  11.620 2.400 11.850 3.720 ;
        RECT  11.360 0.700 11.700 1.465 ;
        RECT  11.395 3.415 11.850 3.720 ;
        END
    END Q
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.625 2.100 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.080 -0.400 12.420 1.005 ;
        RECT  10.470 -0.400 10.810 0.950 ;
        RECT  5.725 -0.400 6.065 0.950 ;
        RECT  0.915 -0.400 1.255 1.395 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  12.080 3.330 12.420 5.280 ;
        RECT  9.800 3.930 10.140 5.280 ;
        RECT  7.185 3.480 7.525 5.280 ;
        RECT  5.885 3.525 6.225 5.280 ;
        RECT  4.585 3.525 4.925 5.280 ;
        RECT  1.940 3.840 2.280 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.645 0.555 0.985 ;
        RECT  0.115 0.645 0.400 2.350 ;
        RECT  0.115 2.120 1.950 2.350 ;
        RECT  1.665 2.120 1.950 2.460 ;
        RECT  0.115 0.645 0.345 3.790 ;
        RECT  0.115 3.450 0.760 3.790 ;
        RECT  2.180 1.090 3.205 1.325 ;
        RECT  0.575 2.855 0.905 3.195 ;
        RECT  0.575 2.930 1.450 3.195 ;
        RECT  1.220 2.930 1.450 4.180 ;
        RECT  2.180 1.090 2.410 3.575 ;
        RECT  1.220 3.345 3.525 3.575 ;
        RECT  3.185 3.345 3.525 3.665 ;
        RECT  1.220 3.345 1.560 4.180 ;
        RECT  1.635 0.630 4.605 0.860 ;
        RECT  4.265 0.630 4.605 1.410 ;
        RECT  1.635 0.630 1.950 1.450 ;
        RECT  6.755 1.240 7.040 2.690 ;
        RECT  6.755 2.460 8.200 2.690 ;
        RECT  7.860 2.460 8.200 2.800 ;
        RECT  2.905 2.290 3.215 3.115 ;
        RECT  6.635 2.720 6.985 3.295 ;
        RECT  2.905 2.885 4.490 3.115 ;
        RECT  6.755 1.240 6.985 3.295 ;
        RECT  4.260 3.065 6.985 3.295 ;
        RECT  6.295 0.780 7.500 1.010 ;
        RECT  4.965 1.070 5.305 1.410 ;
        RECT  6.295 0.780 6.525 1.410 ;
        RECT  4.965 1.180 6.525 1.410 ;
        RECT  2.640 1.555 3.675 1.785 ;
        RECT  7.270 0.780 7.500 2.020 ;
        RECT  2.640 1.555 2.925 1.895 ;
        RECT  7.270 1.790 8.660 2.020 ;
        RECT  7.990 1.790 8.660 2.130 ;
        RECT  3.445 1.555 3.675 2.655 ;
        RECT  6.150 1.180 6.490 2.360 ;
        RECT  3.445 2.290 3.975 2.655 ;
        RECT  6.150 1.180 6.380 2.655 ;
        RECT  3.445 2.425 6.380 2.655 ;
        RECT  5.085 2.425 5.425 2.835 ;
        RECT  8.430 1.790 8.660 3.240 ;
        RECT  8.430 2.900 8.960 3.240 ;
        RECT  7.730 0.630 10.010 0.950 ;
        RECT  7.730 0.630 8.070 0.970 ;
        RECT  8.510 1.220 8.850 1.560 ;
        RECT  8.510 1.330 9.225 1.560 ;
        RECT  8.995 1.330 9.225 2.635 ;
        RECT  8.995 2.405 10.830 2.635 ;
        RECT  10.130 2.405 10.830 2.745 ;
        RECT  10.130 2.405 10.470 3.465 ;
        RECT  9.290 2.405 9.520 3.820 ;
        RECT  8.340 3.480 9.520 3.820 ;
        RECT  9.460 1.180 11.080 1.410 ;
        RECT  10.850 1.180 11.080 1.925 ;
        RECT  11.070 1.695 11.610 1.980 ;
        RECT  9.460 1.180 9.800 2.080 ;
        RECT  11.070 1.695 11.300 3.205 ;
        RECT  10.770 2.975 11.300 3.205 ;
        RECT  10.770 2.975 11.000 4.250 ;
        RECT  10.600 3.930 11.000 4.250 ;
        RECT  1.220 3.345 2.90 3.575 ;
        RECT  1.635 0.630 3.40 0.860 ;
        RECT  4.260 3.065 5.90 3.295 ;
        RECT  3.445 2.425 5.30 2.655 ;
        RECT  7.730 0.630 9.20 0.950 ;
    END
END DFFRQX1

MACRO DFFRQX0
    CLASS CORE ;
    FOREIGN DFFRQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.970 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.577  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.315 2.860 11.845 3.350 ;
        RECT  11.615 0.630 11.845 3.350 ;
        RECT  11.180 0.630 11.845 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.245 4.525 2.630 ;
        END
    END D
    PIN RN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.295  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.500 2.250 10.025 2.815 ;
        END
    END RN
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.215 2.200 5.685 2.630 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.970 5.280 ;
        RECT  11.315 3.810 11.655 5.280 ;
        RECT  9.245 3.910 9.580 5.280 ;
        RECT  6.650 3.630 6.990 5.280 ;
        RECT  4.490 3.910 5.765 5.280 ;
        RECT  0.980 3.520 1.920 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.970 0.400 ;
        RECT  10.380 -0.400 10.720 0.950 ;
        RECT  5.710 -0.400 5.995 1.485 ;
        RECT  0.780 -0.400 1.120 0.980 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 1.970 ;
        RECT  0.115 1.740 2.015 1.970 ;
        RECT  1.730 1.740 2.015 2.460 ;
        RECT  0.115 1.360 0.345 3.860 ;
        RECT  0.115 3.520 0.520 3.860 ;
        RECT  2.245 1.285 3.150 1.590 ;
        RECT  0.630 2.200 0.970 3.060 ;
        RECT  0.630 2.720 2.475 3.060 ;
        RECT  2.245 1.285 2.475 4.250 ;
        RECT  2.245 3.910 3.490 4.250 ;
        RECT  1.580 0.825 4.550 1.055 ;
        RECT  1.580 0.825 1.920 1.510 ;
        RECT  4.210 0.825 4.550 1.545 ;
        RECT  6.685 1.230 6.945 3.200 ;
        RECT  5.865 2.860 7.940 3.200 ;
        RECT  2.870 2.840 3.210 3.675 ;
        RECT  5.865 2.860 6.095 3.675 ;
        RECT  2.870 3.445 6.095 3.675 ;
        RECT  6.225 0.765 7.405 0.995 ;
        RECT  4.825 1.230 5.250 1.945 ;
        RECT  4.825 1.715 6.455 1.945 ;
        RECT  6.225 0.765 6.455 1.950 ;
        RECT  3.445 1.775 4.985 2.005 ;
        RECT  7.175 0.765 7.405 2.530 ;
        RECT  2.705 1.835 3.675 2.180 ;
        RECT  5.990 1.715 6.330 2.395 ;
        RECT  7.175 2.170 8.555 2.530 ;
        RECT  3.445 1.775 3.675 3.180 ;
        RECT  4.755 1.775 4.985 3.200 ;
        RECT  3.445 2.860 3.880 3.180 ;
        RECT  4.755 2.860 5.165 3.200 ;
        RECT  8.270 2.170 8.555 3.450 ;
        RECT  7.635 0.630 9.850 0.860 ;
        RECT  7.635 0.630 7.920 0.970 ;
        RECT  9.510 0.630 9.850 0.970 ;
        RECT  8.480 1.170 8.820 1.510 ;
        RECT  8.785 3.125 10.625 3.465 ;
        RECT  8.785 1.280 9.015 3.970 ;
        RECT  7.950 3.680 9.015 3.970 ;
        RECT  11.065 1.360 11.385 1.920 ;
        RECT  9.430 1.690 11.085 2.020 ;
        RECT  10.855 1.690 11.085 4.250 ;
        RECT  10.065 3.925 11.085 4.250 ;
        RECT  1.580 0.825 3.80 1.055 ;
        RECT  5.865 2.860 6.60 3.200 ;
        RECT  2.870 3.445 5.30 3.675 ;
        RECT  7.635 0.630 8.20 0.860 ;
    END
END DFFRQX0

MACRO DFFQX4
    CLASS CORE ;
    FOREIGN DFFQX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.490 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.221  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.900 2.250 14.365 2.630 ;
        RECT  13.900 2.250 14.240 3.770 ;
        RECT  11.940 2.250 14.365 2.480 ;
        RECT  13.250 1.130 13.590 2.480 ;
        RECT  12.580 2.250 12.920 3.935 ;
        RECT  11.940 1.095 12.170 2.480 ;
        RECT  11.810 1.095 12.170 1.435 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.185  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.240 0.785 2.640 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.505 1.640 5.855 2.100 ;
        RECT  5.165 1.640 5.855 1.970 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 14.490 0.400 ;
        RECT  13.970 -0.400 14.310 1.470 ;
        RECT  12.530 -0.400 12.870 1.470 ;
        RECT  10.310 -0.400 10.650 1.240 ;
        RECT  7.700 -0.400 8.040 1.320 ;
        RECT  5.690 -0.400 6.030 0.950 ;
        RECT  1.580 -0.400 2.400 1.060 ;
        RECT  0.180 -0.400 0.520 0.980 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 14.490 5.280 ;
        RECT  13.340 4.170 13.680 5.280 ;
        RECT  11.820 3.910 12.160 5.280 ;
        RECT  10.555 3.540 10.895 5.280 ;
        RECT  8.460 3.850 8.800 5.280 ;
        RECT  6.040 2.970 6.340 5.280 ;
        RECT  1.995 4.060 2.335 5.280 ;
        RECT  0.940 4.060 1.280 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.375 1.750 2.860 2.090 ;
        RECT  1.375 1.750 1.605 3.370 ;
        RECT  1.375 3.085 1.840 3.370 ;
        RECT  3.090 1.190 3.680 1.530 ;
        RECT  1.835 2.325 3.320 2.665 ;
        RECT  3.090 1.190 3.320 3.275 ;
        RECT  3.090 2.935 3.570 3.275 ;
        RECT  0.180 3.225 0.520 3.830 ;
        RECT  3.950 3.120 4.290 3.830 ;
        RECT  0.180 3.600 4.290 3.830 ;
        RECT  2.630 0.700 4.140 0.930 ;
        RECT  3.910 0.700 4.140 1.550 ;
        RECT  2.630 0.700 2.860 1.520 ;
        RECT  0.780 1.290 2.860 1.520 ;
        RECT  3.910 1.320 4.475 1.550 ;
        RECT  0.780 1.290 1.120 1.630 ;
        RECT  4.155 1.320 4.475 1.660 ;
        RECT  6.320 0.775 7.470 1.005 ;
        RECT  4.370 0.735 5.230 1.075 ;
        RECT  4.705 0.735 5.230 1.410 ;
        RECT  4.705 1.180 6.550 1.410 ;
        RECT  7.240 0.775 7.470 2.090 ;
        RECT  7.240 1.860 8.950 2.090 ;
        RECT  6.320 0.775 6.550 2.100 ;
        RECT  6.235 1.180 6.550 2.100 ;
        RECT  4.705 0.735 4.935 2.430 ;
        RECT  8.610 1.860 8.950 2.200 ;
        RECT  4.705 2.200 5.295 2.430 ;
        RECT  5.065 2.200 5.295 3.195 ;
        RECT  5.065 2.855 5.350 3.195 ;
        RECT  3.635 1.840 3.975 2.180 ;
        RECT  3.635 1.950 4.335 2.180 ;
        RECT  6.780 1.240 7.010 2.860 ;
        RECT  6.780 2.340 7.830 2.680 ;
        RECT  6.780 2.450 9.565 2.680 ;
        RECT  4.105 1.950 4.335 2.890 ;
        RECT  9.280 1.570 9.565 2.680 ;
        RECT  5.580 2.510 7.060 2.740 ;
        RECT  6.720 2.510 7.060 2.860 ;
        RECT  4.105 2.660 4.835 2.890 ;
        RECT  4.570 2.660 4.835 3.655 ;
        RECT  7.930 3.390 9.550 3.620 ;
        RECT  6.720 2.510 6.950 3.855 ;
        RECT  5.580 2.510 5.810 3.655 ;
        RECT  4.570 3.425 5.810 3.655 ;
        RECT  7.930 3.390 8.160 3.855 ;
        RECT  6.720 3.625 8.160 3.855 ;
        RECT  9.210 3.390 9.550 4.000 ;
        RECT  8.850 0.920 9.190 1.340 ;
        RECT  8.850 1.110 10.025 1.340 ;
        RECT  10.910 2.120 11.250 2.460 ;
        RECT  9.795 2.230 11.250 2.460 ;
        RECT  7.380 2.930 10.025 3.160 ;
        RECT  7.270 3.110 7.610 3.395 ;
        RECT  9.795 1.110 10.025 3.880 ;
        RECT  9.780 2.930 10.025 3.880 ;
        RECT  9.780 3.540 10.120 3.880 ;
        RECT  11.110 0.900 11.450 1.890 ;
        RECT  10.255 1.550 11.450 1.890 ;
        RECT  10.255 1.660 11.710 1.890 ;
        RECT  11.480 1.660 11.710 3.510 ;
        RECT  11.260 2.690 11.710 3.510 ;
        RECT  0.180 3.600 3.50 3.830 ;
        RECT  0.780 1.290 1.00 1.520 ;
        RECT  6.780 2.450 8.40 2.680 ;
        RECT  7.380 2.930 9.60 3.160 ;
    END
END DFFQX4

MACRO DFFQX2
    CLASS CORE ;
    FOREIGN DFFQX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.205 1.240 10.600 3.550 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.635 3.770 2.115 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 1.640 4.915 2.180 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.820 3.950 11.160 5.280 ;
        RECT  9.500 3.495 9.840 5.280 ;
        RECT  8.295 3.490 8.635 5.280 ;
        RECT  5.910 3.830 6.250 5.280 ;
        RECT  4.770 3.910 5.110 5.280 ;
        RECT  3.510 3.880 3.850 5.280 ;
        RECT  1.680 3.960 2.020 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.820 -0.400 11.160 0.720 ;
        RECT  9.700 -0.400 10.040 0.720 ;
        RECT  8.300 -0.400 8.640 1.060 ;
        RECT  6.650 -0.400 6.990 0.950 ;
        RECT  4.640 -0.400 4.975 0.950 ;
        RECT  3.080 -0.400 3.420 0.840 ;
        RECT  0.700 -0.400 1.040 1.010 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.360 0.520 2.870 ;
        RECT  0.115 2.640 1.455 2.870 ;
        RECT  1.115 2.640 1.455 2.925 ;
        RECT  0.115 1.360 0.345 3.940 ;
        RECT  0.115 3.710 1.280 3.940 ;
        RECT  0.940 3.710 1.280 4.070 ;
        RECT  1.270 0.630 2.350 0.950 ;
        RECT  1.270 0.630 1.500 2.410 ;
        RECT  1.270 2.180 1.675 2.410 ;
        RECT  1.625 2.185 1.915 2.415 ;
        RECT  0.575 3.100 0.860 3.440 ;
        RECT  1.685 2.185 1.915 3.625 ;
        RECT  0.575 3.210 1.915 3.440 ;
        RECT  1.685 3.395 2.820 3.625 ;
        RECT  2.480 3.395 2.820 3.735 ;
        RECT  5.665 1.195 5.950 1.870 ;
        RECT  5.775 2.560 6.925 2.900 ;
        RECT  2.145 2.360 2.430 3.165 ;
        RECT  2.145 2.935 3.700 3.165 ;
        RECT  3.470 2.935 3.700 3.410 ;
        RECT  5.530 2.860 6.005 3.410 ;
        RECT  5.775 1.695 6.005 3.410 ;
        RECT  3.470 3.180 6.005 3.410 ;
        RECT  5.205 0.735 6.420 0.965 ;
        RECT  6.190 0.735 6.420 1.555 ;
        RECT  3.880 1.180 5.435 1.410 ;
        RECT  3.880 1.090 4.220 1.430 ;
        RECT  6.190 1.325 7.350 1.555 ;
        RECT  1.730 1.670 2.990 1.955 ;
        RECT  5.205 0.735 5.435 2.420 ;
        RECT  5.175 1.180 5.435 2.420 ;
        RECT  7.120 1.325 7.350 2.190 ;
        RECT  2.760 1.670 2.990 2.705 ;
        RECT  5.175 2.080 5.500 2.420 ;
        RECT  2.760 2.340 3.100 2.705 ;
        RECT  4.000 1.180 4.230 2.950 ;
        RECT  2.760 2.475 4.230 2.705 ;
        RECT  4.000 2.610 4.550 2.950 ;
        RECT  7.265 1.850 7.550 3.310 ;
        RECT  7.475 0.720 8.010 1.060 ;
        RECT  8.920 2.120 9.260 2.460 ;
        RECT  7.780 2.230 9.260 2.460 ;
        RECT  7.780 0.720 8.010 4.005 ;
        RECT  7.065 3.665 8.010 4.005 ;
        RECT  9.000 0.650 9.340 1.180 ;
        RECT  9.000 0.950 9.720 1.180 ;
        RECT  9.490 0.950 9.720 2.960 ;
        RECT  8.240 2.730 9.720 2.960 ;
        RECT  8.240 2.730 9.280 3.070 ;
        RECT  3.470 3.180 5.50 3.410 ;
    END
END DFFQX2

MACRO DFFQX1
    CLASS CORE ;
    FOREIGN DFFQX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.189  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.070 1.030 3.395 2.010 ;
        RECT  2.645 1.030 3.395 1.410 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.662  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.640 2.400 10.585 2.630 ;
        RECT  9.970 2.250 10.585 2.630 ;
        RECT  9.970 1.320 10.200 2.630 ;
        RECT  9.380 1.320 10.200 1.550 ;
        RECT  9.380 3.325 9.870 3.610 ;
        RECT  9.640 2.400 9.870 3.610 ;
        RECT  9.380 0.700 9.720 1.550 ;
        END
    END Q
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.297  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.340 2.140 ;
        END
    END CN
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  10.100 -0.400 10.440 1.090 ;
        RECT  8.575 -0.400 8.915 1.440 ;
        RECT  6.995 -0.400 7.335 0.790 ;
        RECT  4.520 -0.400 4.860 0.925 ;
        RECT  3.060 -0.400 3.400 0.800 ;
        RECT  0.960 -0.400 1.300 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.100 3.330 10.440 5.280 ;
        RECT  8.040 4.145 8.380 5.280 ;
        RECT  5.820 3.810 6.160 5.280 ;
        RECT  4.690 3.525 5.030 5.280 ;
        RECT  3.590 3.810 3.930 5.280 ;
        RECT  1.220 4.170 1.560 5.280 ;
        RECT  0.420 4.170 0.760 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.115 0.645 0.520 2.480 ;
        RECT  0.115 2.140 1.020 2.480 ;
        RECT  0.115 0.645 0.345 3.790 ;
        RECT  0.115 3.450 0.760 3.790 ;
        RECT  1.860 0.630 2.200 1.410 ;
        RECT  1.250 1.180 2.200 1.410 ;
        RECT  0.700 2.880 1.480 3.220 ;
        RECT  1.250 1.180 1.480 3.875 ;
        RECT  1.250 3.645 2.530 3.875 ;
        RECT  2.190 3.645 2.530 3.985 ;
        RECT  5.550 1.240 5.835 1.580 ;
        RECT  5.605 1.240 5.835 2.800 ;
        RECT  5.605 2.460 6.870 2.800 ;
        RECT  1.970 2.565 2.310 3.360 ;
        RECT  5.450 2.540 5.810 3.295 ;
        RECT  3.575 3.065 5.810 3.295 ;
        RECT  1.970 3.130 3.755 3.360 ;
        RECT  5.090 0.780 6.295 1.010 ;
        RECT  3.760 1.070 4.100 1.385 ;
        RECT  5.090 0.780 5.320 1.385 ;
        RECT  3.760 1.155 5.320 1.385 ;
        RECT  6.065 0.780 6.295 1.905 ;
        RECT  1.710 1.685 2.050 2.025 ;
        RECT  6.065 1.675 7.130 1.905 ;
        RECT  6.785 1.765 7.505 2.015 ;
        RECT  1.710 1.795 2.840 2.025 ;
        RECT  4.945 1.155 5.290 2.310 ;
        RECT  2.610 1.795 2.840 2.900 ;
        RECT  4.945 1.155 5.175 2.765 ;
        RECT  2.610 2.535 5.175 2.765 ;
        RECT  3.890 2.535 4.230 2.835 ;
        RECT  7.275 1.765 7.505 3.240 ;
        RECT  2.610 2.535 2.980 2.900 ;
        RECT  7.275 2.900 7.630 3.240 ;
        RECT  7.305 1.150 7.645 1.490 ;
        RECT  7.305 1.260 7.965 1.490 ;
        RECT  7.735 1.260 7.965 2.580 ;
        RECT  7.860 2.350 8.940 2.635 ;
        RECT  7.860 2.350 8.090 3.785 ;
        RECT  7.010 3.555 8.090 3.785 ;
        RECT  7.010 3.555 7.350 3.895 ;
        RECT  8.255 1.670 8.595 2.010 ;
        RECT  8.255 1.780 9.720 2.010 ;
        RECT  9.180 1.780 9.720 2.120 ;
        RECT  9.180 1.780 9.410 3.095 ;
        RECT  8.840 2.865 9.410 3.095 ;
        RECT  8.840 2.865 9.150 4.200 ;
        RECT  8.840 3.860 9.180 4.200 ;
        RECT  3.575 3.065 4.10 3.295 ;
        RECT  2.610 2.535 4.40 2.765 ;
    END
END DFFQX1

MACRO DFFQX0
    CLASS CORE ;
    FOREIGN DFFQX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.493  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.520 2.250 9.955 3.085 ;
        RECT  9.725 0.630 9.955 3.085 ;
        RECT  9.030 0.630 9.955 0.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.130 2.220 3.655 2.685 ;
        END
    END D
    PIN CN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.345 2.160 4.865 2.640 ;
        END
    END CN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  9.445 3.545 9.785 5.280 ;
        RECT  8.055 3.880 8.395 5.280 ;
        RECT  5.300 3.650 5.640 5.280 ;
        RECT  3.490 3.910 4.760 5.280 ;
        RECT  0.780 4.075 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.190 -0.400 8.570 0.970 ;
        RECT  6.510 -0.400 6.795 0.970 ;
        RECT  4.560 -0.400 4.845 0.970 ;
        RECT  3.260 -0.400 3.600 0.970 ;
        RECT  0.780 -0.400 1.120 0.940 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.115 1.255 0.520 2.420 ;
        RECT  0.115 2.040 1.275 2.420 ;
        RECT  0.115 1.255 0.345 3.700 ;
        RECT  0.115 3.360 0.520 3.700 ;
        RECT  1.505 1.165 2.540 1.505 ;
        RECT  1.505 1.165 1.735 2.805 ;
        RECT  0.575 2.790 1.640 3.130 ;
        RECT  1.410 2.615 1.640 4.120 ;
        RECT  1.410 3.890 2.360 4.120 ;
        RECT  2.020 3.890 2.360 4.230 ;
        RECT  5.555 1.270 5.820 1.905 ;
        RECT  5.675 1.675 5.905 3.200 ;
        RECT  5.285 2.860 6.635 3.200 ;
        RECT  4.455 2.945 6.635 3.200 ;
        RECT  1.870 3.020 2.210 3.360 ;
        RECT  1.980 3.020 2.210 3.660 ;
        RECT  4.455 2.945 4.685 3.660 ;
        RECT  1.980 3.430 4.685 3.660 ;
        RECT  5.075 0.810 6.280 1.040 ;
        RECT  3.885 1.270 4.300 1.610 ;
        RECT  6.050 0.810 6.280 1.445 ;
        RECT  5.075 0.810 5.325 1.610 ;
        RECT  3.885 1.380 5.325 1.610 ;
        RECT  1.965 1.735 4.115 1.965 ;
        RECT  1.965 1.735 2.770 2.105 ;
        RECT  6.235 1.215 6.465 2.530 ;
        RECT  5.095 0.810 5.325 2.575 ;
        RECT  6.235 2.190 6.590 2.530 ;
        RECT  6.235 2.230 7.245 2.530 ;
        RECT  5.095 2.220 5.445 2.575 ;
        RECT  2.540 1.735 2.770 3.180 ;
        RECT  3.885 1.270 4.115 3.200 ;
        RECT  7.015 2.230 7.245 3.445 ;
        RECT  2.540 2.840 2.880 3.180 ;
        RECT  3.820 2.860 4.160 3.200 ;
        RECT  7.015 3.105 7.365 3.445 ;
        RECT  7.330 0.630 7.825 0.970 ;
        RECT  7.595 2.570 8.830 2.800 ;
        RECT  8.490 2.570 8.830 2.910 ;
        RECT  7.595 0.630 7.825 3.990 ;
        RECT  6.700 3.675 7.825 3.990 ;
        RECT  9.010 1.360 9.370 1.700 ;
        RECT  9.010 1.360 9.290 2.130 ;
        RECT  8.080 1.900 9.290 2.130 ;
        RECT  8.080 1.900 8.420 2.240 ;
        RECT  9.060 1.360 9.290 3.370 ;
        RECT  8.555 3.140 9.290 3.370 ;
        RECT  8.555 3.140 8.895 3.480 ;
        RECT  4.455 2.945 5.60 3.200 ;
        RECT  1.980 3.430 3.40 3.660 ;
        RECT  1.965 1.735 3.80 1.965 ;
    END
END DFFQX0

MACRO DECAP7LP
    CLASS CORE SPACER ;
    FOREIGN DECAP7LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.280 -0.400 3.620 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  0.790 2.740 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.775 1.305 1.130 2.510 ;
        RECT  3.280 1.825 3.635 3.910 ;
    END
END DECAP7LP

MACRO DECAP7
    CLASS CORE SPACER ;
    FOREIGN DECAP7 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.890 -0.400 4.230 1.510 ;
        RECT  0.940 -0.400 1.280 1.510 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.130 3.370 3.470 5.280 ;
        RECT  0.180 3.370 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.795 0.520 2.555 ;
        RECT  0.165 2.215 0.975 2.555 ;
        RECT  3.435 1.785 4.245 2.125 ;
        RECT  3.890 1.785 4.245 3.545 ;
    END
END DECAP7

MACRO DECAP5LP
    CLASS CORE SPACER ;
    FOREIGN DECAP5LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.020 -0.400 2.360 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.790 2.740 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.775 1.305 1.130 2.510 ;
        RECT  2.020 1.825 2.375 3.910 ;
    END
END DECAP5LP

MACRO DECAP5
    CLASS CORE SPACER ;
    FOREIGN DECAP5 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 1.180 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.180 3.700 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.810 0.520 2.510 ;
        RECT  0.165 2.170 0.975 2.510 ;
        RECT  2.175 1.800 2.985 2.140 ;
        RECT  2.630 1.800 2.985 3.565 ;
    END
END DECAP5

MACRO DECAP3
    CLASS CORE SPACER ;
    FOREIGN DECAP3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.890 0.400 ;
        RECT  1.370 -0.400 1.710 1.180 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.890 5.280 ;
        RECT  0.180 3.700 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.835 0.520 2.510 ;
        RECT  1.370 1.825 1.725 3.555 ;
    END
END DECAP3

MACRO DECAP25LP
    CLASS CORE SPACER ;
    FOREIGN DECAP25LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  14.620 -0.400 14.960 1.310 ;
        RECT  12.465 -0.400 12.805 1.310 ;
        RECT  10.310 -0.400 10.650 1.310 ;
        RECT  8.155 -0.400 8.495 1.310 ;
        RECT  6.000 -0.400 6.340 1.310 ;
        RECT  3.835 -0.400 4.175 1.310 ;
        RECT  1.680 -0.400 2.020 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  13.730 3.570 14.070 5.280 ;
        RECT  11.565 3.570 11.905 5.280 ;
        RECT  9.410 3.570 9.750 5.280 ;
        RECT  7.255 3.570 7.595 5.280 ;
        RECT  5.100 3.570 5.440 5.280 ;
        RECT  2.945 3.570 3.285 5.280 ;
        RECT  0.790 3.570 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.775 1.265 1.130 2.555 ;
        RECT  0.775 2.215 1.585 2.555 ;
        RECT  14.165 1.785 14.975 2.125 ;
        RECT  14.620 1.785 14.975 3.075 ;
    END
END DECAP25LP

MACRO DECAP25
    CLASS CORE SPACER ;
    FOREIGN DECAP25 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        RECT  15.230 -0.400 15.570 1.510 ;
        RECT  12.845 -0.400 13.185 1.510 ;
        RECT  10.465 -0.400 10.805 1.510 ;
        RECT  8.080 -0.400 8.420 1.510 ;
        RECT  5.700 -0.400 6.040 1.510 ;
        RECT  3.320 -0.400 3.660 1.510 ;
        RECT  0.940 -0.400 1.280 1.510 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        RECT  14.470 3.370 14.810 5.280 ;
        RECT  12.080 3.370 12.420 5.280 ;
        RECT  9.700 3.370 10.040 5.280 ;
        RECT  7.320 3.370 7.660 5.280 ;
        RECT  4.940 3.370 5.280 5.280 ;
        RECT  2.560 3.370 2.900 5.280 ;
        RECT  0.180 3.370 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.795 0.520 2.555 ;
        RECT  0.165 2.215 0.975 2.555 ;
        RECT  14.775 1.785 15.585 2.125 ;
        RECT  15.230 1.785 15.585 3.545 ;
    END
END DECAP25

MACRO DECAP15LP
    CLASS CORE SPACER ;
    FOREIGN DECAP15LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.320 -0.400 8.660 1.310 ;
        RECT  6.110 -0.400 6.450 1.310 ;
        RECT  3.890 -0.400 4.230 1.310 ;
        RECT  1.680 -0.400 2.020 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  7.430 3.570 7.770 5.280 ;
        RECT  5.220 3.570 5.560 5.280 ;
        RECT  3.000 3.570 3.340 5.280 ;
        RECT  0.790 3.570 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.775 1.265 1.130 2.555 ;
        RECT  0.775 2.215 1.585 2.555 ;
        RECT  7.865 1.785 8.675 2.125 ;
        RECT  8.320 1.785 8.675 3.075 ;
    END
END DECAP15LP

MACRO DECAP15
    CLASS CORE SPACER ;
    FOREIGN DECAP15 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.930 -0.400 9.270 1.510 ;
        RECT  6.260 -0.400 6.600 1.510 ;
        RECT  3.600 -0.400 3.940 1.510 ;
        RECT  0.940 -0.400 1.280 1.510 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.170 3.370 8.510 5.280 ;
        RECT  5.510 3.370 5.850 5.280 ;
        RECT  2.850 3.370 3.190 5.280 ;
        RECT  0.180 3.370 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.795 0.520 2.555 ;
        RECT  0.165 2.215 0.975 2.555 ;
        RECT  8.475 1.785 9.285 2.125 ;
        RECT  8.930 1.785 9.285 3.545 ;
    END
END DECAP15

MACRO DECAP10LP
    CLASS CORE SPACER ;
    FOREIGN DECAP10LP 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.170 -0.400 5.510 1.310 ;
        RECT  1.680 -0.400 2.020 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  4.280 3.570 4.620 5.280 ;
        RECT  0.790 3.570 1.130 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.775 1.265 1.130 2.555 ;
        RECT  0.775 2.215 1.585 2.555 ;
        RECT  4.715 1.785 5.525 2.125 ;
        RECT  5.170 1.785 5.525 3.075 ;
    END
END DECAP10LP

MACRO DECAP10
    CLASS CORE SPACER ;
    FOREIGN DECAP10 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 1.510 ;
        RECT  3.360 -0.400 3.700 1.510 ;
        RECT  0.940 -0.400 1.280 1.510 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.020 3.370 5.360 5.280 ;
        RECT  2.600 3.370 2.940 5.280 ;
        RECT  0.180 3.370 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.165 0.795 0.520 2.555 ;
        RECT  0.165 2.215 0.975 2.555 ;
        RECT  5.325 1.785 6.135 2.125 ;
        RECT  5.780 1.785 6.135 3.545 ;
    END
END DECAP10

MACRO BUX8
    CLASS CORE ;
    FOREIGN BUX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.518  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.300 0.905 8.640 4.180 ;
        RECT  5.380 1.560 8.640 2.060 ;
        RECT  6.820 0.905 7.165 2.060 ;
        RECT  6.820 0.905 7.160 4.180 ;
        RECT  5.380 0.905 5.720 4.180 ;
        RECT  3.940 2.365 5.720 2.705 ;
        RECT  3.940 1.270 5.720 1.560 ;
        RECT  3.940 2.365 4.280 4.180 ;
        RECT  3.940 0.905 4.280 1.560 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.696  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.555 0.550 2.365 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.540 -0.400 7.880 1.245 ;
        RECT  6.100 -0.400 6.440 1.245 ;
        RECT  4.660 -0.400 5.000 1.040 ;
        RECT  3.135 -0.400 3.475 1.245 ;
        RECT  1.650 -0.400 1.995 1.245 ;
        RECT  0.210 -0.400 0.550 1.245 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.540 2.315 7.880 5.280 ;
        RECT  6.100 2.315 6.440 5.280 ;
        RECT  4.660 2.935 5.000 5.280 ;
        RECT  3.160 2.660 3.500 5.280 ;
        RECT  1.650 2.660 2.000 5.280 ;
        RECT  0.210 2.660 0.550 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.930 1.795 5.035 2.135 ;
        RECT  0.930 0.905 1.270 4.180 ;
        RECT  2.370 0.905 2.710 4.180 ;
        RECT  0.930 1.795 4.40 2.135 ;
    END
END BUX8

MACRO BUX6
    CLASS CORE ;
    FOREIGN BUX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.054  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 0.905 6.750 4.180 ;
        RECT  3.570 1.560 6.750 2.060 ;
        RECT  4.930 0.905 5.275 2.060 ;
        RECT  4.930 0.905 5.270 4.180 ;
        RECT  3.490 2.310 3.830 4.180 ;
        RECT  3.570 0.905 3.830 4.180 ;
        RECT  3.490 0.905 3.830 1.245 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.520 1.325 2.020 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.650 -0.400 5.990 1.245 ;
        RECT  4.210 -0.400 4.550 1.245 ;
        RECT  2.565 -0.400 2.910 1.320 ;
        RECT  0.900 -0.400 1.245 1.245 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.650 2.310 5.990 5.280 ;
        RECT  4.210 2.310 4.550 5.280 ;
        RECT  2.340 2.670 3.110 5.280 ;
        RECT  2.770 2.310 3.110 5.280 ;
        RECT  0.900 2.780 1.250 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.620 1.705 3.340 2.045 ;
        RECT  0.180 2.250 1.960 2.530 ;
        RECT  0.180 0.905 0.520 4.180 ;
        RECT  1.620 0.905 1.960 4.180 ;
    END
END BUX6

MACRO BUX4
    CLASS CORE ;
    FOREIGN BUX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.441  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.800 0.905 4.145 4.160 ;
        RECT  2.415 1.600 4.145 2.060 ;
        RECT  2.360 2.640 2.700 4.160 ;
        RECT  2.415 0.905 2.700 4.160 ;
        RECT  2.360 0.905 2.700 1.245 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.846  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.505 0.550 2.065 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.520 -0.400 4.860 1.245 ;
        RECT  3.080 -0.400 3.420 1.245 ;
        RECT  1.635 -0.400 1.980 1.245 ;
        RECT  0.200 -0.400 0.545 1.245 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.520 2.635 4.860 5.280 ;
        RECT  3.080 2.635 3.420 5.280 ;
        RECT  1.640 2.640 1.980 5.280 ;
        RECT  0.200 2.640 0.540 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.920 1.550 2.170 2.360 ;
        RECT  0.920 0.905 1.260 4.160 ;
    END
END BUX4

MACRO BUX3
    CLASS CORE ;
    FOREIGN BUX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 0.975 4.235 4.160 ;
        RECT  2.505 1.600 4.235 2.060 ;
        RECT  2.450 2.640 2.790 4.160 ;
        RECT  2.505 0.975 2.790 4.160 ;
        RECT  2.450 0.975 2.790 1.315 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.637  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.505 0.550 2.065 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.170 -0.400 3.510 1.315 ;
        RECT  1.730 -0.400 2.070 1.315 ;
        RECT  0.290 -0.400 0.635 1.250 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.170 2.635 3.510 5.280 ;
        RECT  1.730 2.640 2.070 5.280 ;
        RECT  0.290 2.640 0.630 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.010 1.550 2.260 2.360 ;
        RECT  1.010 0.910 1.350 3.760 ;
    END
END BUX3

MACRO BUX20
    CLASS CORE ;
    FOREIGN BUX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 4.230  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.790 2.140 2.130 ;
        RECT  0.125 1.640 0.505 2.130 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.715  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  19.640 0.905 19.980 4.160 ;
        RECT  12.420 1.510 19.980 2.310 ;
        RECT  18.180 0.905 18.520 4.160 ;
        RECT  16.740 0.920 17.080 4.140 ;
        RECT  15.300 0.920 15.640 4.160 ;
        RECT  13.860 0.920 14.200 4.160 ;
        RECT  12.420 0.920 12.760 4.160 ;
        RECT  8.100 2.375 12.760 2.715 ;
        RECT  8.100 1.285 12.760 1.575 ;
        RECT  10.980 2.375 11.320 4.160 ;
        RECT  10.980 0.920 11.320 1.575 ;
        RECT  9.540 0.920 9.885 1.575 ;
        RECT  9.540 2.375 9.880 4.160 ;
        RECT  8.100 2.375 8.440 4.160 ;
        RECT  8.100 0.920 8.440 1.575 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 20.160 0.400 ;
        RECT  18.900 -0.400 19.240 1.245 ;
        RECT  17.460 -0.400 17.800 1.260 ;
        RECT  16.020 -0.400 16.360 1.260 ;
        RECT  14.580 -0.400 14.920 1.260 ;
        RECT  13.140 -0.400 13.480 1.260 ;
        RECT  11.700 -0.400 12.040 1.055 ;
        RECT  10.260 -0.400 10.600 1.055 ;
        RECT  8.820 -0.400 10.600 0.405 ;
        RECT  8.820 -0.400 9.160 1.055 ;
        RECT  7.380 -0.400 7.720 1.390 ;
        RECT  5.940 -0.400 6.280 1.260 ;
        RECT  4.500 -0.400 4.840 1.260 ;
        RECT  3.060 -0.400 3.400 1.250 ;
        RECT  1.615 -0.400 1.960 1.060 ;
        RECT  0.180 -0.400 0.520 1.260 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 20.160 5.280 ;
        RECT  18.900 2.620 19.240 5.280 ;
        RECT  17.460 2.540 17.800 5.280 ;
        RECT  16.020 2.560 16.360 5.280 ;
        RECT  14.580 2.560 14.920 5.280 ;
        RECT  13.140 2.560 13.480 5.280 ;
        RECT  11.700 2.945 12.040 5.280 ;
        RECT  10.260 2.945 10.600 5.280 ;
        RECT  8.820 2.945 9.160 5.280 ;
        RECT  7.380 2.640 7.730 5.280 ;
        RECT  5.940 2.640 6.280 5.280 ;
        RECT  4.500 2.640 4.840 5.280 ;
        RECT  3.060 2.640 3.400 5.280 ;
        RECT  1.620 2.875 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 0.920 1.240 1.560 ;
        RECT  2.340 0.920 2.680 1.560 ;
        RECT  0.900 1.290 2.680 1.560 ;
        RECT  2.370 1.805 12.190 2.145 ;
        RECT  0.900 2.360 2.680 2.645 ;
        RECT  0.900 2.360 1.240 4.160 ;
        RECT  2.370 0.920 2.680 4.160 ;
        RECT  2.340 2.360 2.680 4.160 ;
        RECT  3.780 0.920 4.120 4.160 ;
        RECT  5.220 0.920 5.560 4.160 ;
        RECT  6.660 0.920 7.000 4.160 ;
        RECT  2.370 1.805 11.40 2.145 ;
    END
END BUX20

MACRO BUX2
    CLASS CORE ;
    FOREIGN BUX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.423  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.640 0.505 2.225 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.220  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.920 1.640 2.395 2.020 ;
        RECT  1.910 2.660 2.250 4.180 ;
        RECT  1.920 0.905 2.250 4.180 ;
        RECT  1.910 0.905 2.250 1.245 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 1.245 ;
        RECT  1.190 -0.400 1.530 1.130 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  2.630 2.655 2.970 5.280 ;
        RECT  1.190 2.735 1.530 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.430 0.905 0.770 1.410 ;
        RECT  0.735 1.720 1.690 2.060 ;
        RECT  0.735 1.180 0.965 2.685 ;
        RECT  0.430 2.455 0.770 4.180 ;
    END
END BUX2

MACRO BUX16
    CLASS CORE ;
    FOREIGN BUX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.384  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.805 1.915 2.145 ;
        RECT  0.125 1.640 0.505 2.145 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.025  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.730 0.920 16.070 4.160 ;
        RECT  9.850 1.440 16.070 2.140 ;
        RECT  14.250 0.920 14.595 2.140 ;
        RECT  14.250 0.920 14.590 4.160 ;
        RECT  12.770 0.920 13.110 4.160 ;
        RECT  11.290 0.920 11.635 2.140 ;
        RECT  11.290 0.920 11.630 4.160 ;
        RECT  9.850 0.920 10.190 4.160 ;
        RECT  6.930 2.390 10.190 2.730 ;
        RECT  6.930 1.285 10.190 1.590 ;
        RECT  8.370 0.920 8.715 1.590 ;
        RECT  8.370 2.390 8.710 4.160 ;
        RECT  6.930 2.390 7.270 4.160 ;
        RECT  6.930 0.920 7.270 1.590 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  16.490 -0.400 16.830 1.260 ;
        RECT  14.970 -0.400 15.310 1.190 ;
        RECT  13.530 -0.400 13.870 1.190 ;
        RECT  12.010 -0.400 12.350 1.190 ;
        RECT  10.570 -0.400 10.910 1.190 ;
        RECT  9.090 -0.400 9.430 1.055 ;
        RECT  7.650 -0.400 7.990 1.055 ;
        RECT  6.090 -0.400 6.430 1.260 ;
        RECT  4.500 -0.400 4.845 1.260 ;
        RECT  3.060 -0.400 3.405 1.260 ;
        RECT  1.615 -0.400 1.960 1.055 ;
        RECT  0.175 -0.400 0.520 1.260 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  16.490 2.760 16.845 5.280 ;
        RECT  14.970 2.390 15.310 5.280 ;
        RECT  13.530 2.390 13.870 5.280 ;
        RECT  12.010 2.390 12.350 5.280 ;
        RECT  10.570 2.390 10.910 5.280 ;
        RECT  9.090 2.960 9.430 5.280 ;
        RECT  7.650 2.960 7.990 5.280 ;
        RECT  6.095 2.390 6.440 5.280 ;
        RECT  4.500 2.640 4.840 5.280 ;
        RECT  3.060 2.640 3.400 5.280 ;
        RECT  1.620 2.880 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.895 0.920 1.240 1.575 ;
        RECT  0.895 1.285 2.680 1.575 ;
        RECT  2.335 1.820 9.600 2.160 ;
        RECT  0.895 2.375 2.680 2.650 ;
        RECT  0.895 2.375 1.240 4.160 ;
        RECT  2.335 0.920 2.680 4.160 ;
        RECT  3.775 0.920 4.120 4.160 ;
        RECT  5.215 0.920 5.560 4.160 ;
        RECT  2.335 1.820 8.30 2.160 ;
    END
END BUX16

MACRO BUX12
    CLASS CORE ;
    FOREIGN BUX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.312  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  11.320 0.905 11.660 4.180 ;
        RECT  8.400 1.500 11.660 2.100 ;
        RECT  9.840 0.905 10.185 2.100 ;
        RECT  9.840 0.905 10.180 4.180 ;
        RECT  8.400 0.905 8.740 4.180 ;
        RECT  5.480 2.360 8.740 2.650 ;
        RECT  5.480 1.270 8.740 1.560 ;
        RECT  6.920 0.905 7.265 1.560 ;
        RECT  6.920 2.360 7.260 4.180 ;
        RECT  5.480 0.905 5.825 1.560 ;
        RECT  5.480 2.360 5.820 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.538  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.520 0.550 2.360 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.080 -0.400 12.420 1.245 ;
        RECT  10.560 -0.400 10.900 1.245 ;
        RECT  9.120 -0.400 9.460 1.245 ;
        RECT  7.640 -0.400 7.980 1.040 ;
        RECT  6.200 -0.400 6.540 1.040 ;
        RECT  4.640 -0.400 4.980 1.245 ;
        RECT  3.060 -0.400 3.405 1.245 ;
        RECT  1.615 -0.400 1.960 1.245 ;
        RECT  0.175 -0.400 0.520 1.245 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  12.080 2.760 12.435 5.280 ;
        RECT  10.560 2.330 10.900 5.280 ;
        RECT  9.120 2.330 9.460 5.280 ;
        RECT  7.640 2.880 7.980 5.280 ;
        RECT  6.200 2.880 6.540 5.280 ;
        RECT  4.645 2.360 4.990 5.280 ;
        RECT  3.060 2.660 3.410 5.280 ;
        RECT  1.610 2.660 1.960 5.280 ;
        RECT  0.180 2.660 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.790 8.170 2.130 ;
        RECT  0.900 0.905 1.240 4.180 ;
        RECT  2.340 0.905 2.680 4.180 ;
        RECT  3.780 0.905 4.120 4.180 ;
        RECT  0.900 1.790 7.20 2.130 ;
    END
END BUX12

MACRO BUX1
    CLASS CORE ;
    FOREIGN BUX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.085  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.735 1.640 2.395 2.020 ;
        RECT  1.700 2.640 2.045 4.160 ;
        RECT  1.735 1.050 2.045 4.160 ;
        RECT  1.700 1.050 2.045 1.390 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.212  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 3.460 0.750 3.880 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.975 -0.400 1.320 1.390 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.980 2.635 1.320 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.810 1.480 2.150 ;
        RECT  0.180 1.170 0.520 3.170 ;
    END
END BUX1

MACRO BUX0
    CLASS CORE ;
    FOREIGN BUX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.621  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.835 2.250 2.395 2.630 ;
        RECT  1.780 2.640 2.120 2.980 ;
        RECT  1.835 1.170 2.120 2.980 ;
        RECT  1.780 1.170 2.120 1.510 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 3.465 0.750 3.855 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.980 2.745 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.975 -0.400 1.320 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.810 1.590 2.150 ;
        RECT  0.180 1.170 0.520 2.980 ;
    END
END BUX0

MACRO BUCX8
    CLASS CORE ;
    FOREIGN BUCX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.073  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.950 0.700 7.435 4.180 ;
        RECT  4.070 1.740 7.435 2.240 ;
        RECT  5.500 1.740 5.870 4.180 ;
        RECT  5.510 0.700 5.850 4.180 ;
        RECT  4.070 0.915 4.410 4.180 ;
        RECT  2.630 3.100 4.410 3.380 ;
        RECT  2.630 3.100 2.970 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.894  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.600 2.460 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 1.510 ;
        RECT  6.230 -0.400 6.570 1.510 ;
        RECT  4.790 -0.400 5.130 1.510 ;
        RECT  3.350 -0.400 3.690 1.190 ;
        RECT  1.380 -0.400 1.720 1.510 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.670 2.640 8.010 5.280 ;
        RECT  6.230 2.490 6.570 5.280 ;
        RECT  4.790 2.490 5.130 5.280 ;
        RECT  3.340 3.610 3.690 5.280 ;
        RECT  0.180 3.960 2.170 5.280 ;
        RECT  1.830 3.490 2.170 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.480 1.040 1.150 1.380 ;
        RECT  0.850 1.930 3.265 2.270 ;
        RECT  0.850 1.040 1.150 3.560 ;
        RECT  0.740 2.645 1.150 3.560 ;
        RECT  2.260 0.630 3.120 1.700 ;
        RECT  2.260 1.420 3.775 1.700 ;
        RECT  3.495 1.420 3.775 2.780 ;
        RECT  2.070 2.500 3.775 2.780 ;
        RECT  2.070 2.500 2.410 2.990 ;
        RECT  0.850 1.930 2.80 2.270 ;
    END
END BUCX8

MACRO BUCX6
    CLASS CORE ;
    FOREIGN BUCX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.851  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.600 0.760 2.410 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.694  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.680 1.810 6.175 4.180 ;
        RECT  5.690 0.700 6.175 4.180 ;
        RECT  4.250 1.810 6.175 2.310 ;
        RECT  4.250 0.700 4.590 4.180 ;
        RECT  2.810 3.020 4.590 3.320 ;
        RECT  2.810 3.020 3.150 4.180 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 1.325 ;
        RECT  4.970 -0.400 5.310 1.510 ;
        RECT  3.530 -0.400 3.870 1.040 ;
        RECT  1.530 -0.400 1.870 1.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 2.640 6.750 5.280 ;
        RECT  4.970 2.550 5.310 5.280 ;
        RECT  3.530 3.550 3.870 5.280 ;
        RECT  1.610 3.120 2.430 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.600 1.015 1.300 1.355 ;
        RECT  1.010 1.810 3.440 2.150 ;
        RECT  1.010 1.015 1.300 3.460 ;
        RECT  0.900 2.640 1.300 3.460 ;
        RECT  2.440 0.860 3.300 1.200 ;
        RECT  2.960 0.630 3.300 1.520 ;
        RECT  2.960 1.270 3.970 1.520 ;
        RECT  3.670 1.270 3.970 2.720 ;
        RECT  2.270 2.380 3.970 2.720 ;
        RECT  1.010 1.810 2.80 2.150 ;
    END
END BUCX6

MACRO BUCX4
    CLASS CORE ;
    FOREIGN BUCX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.726  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.760 2.075 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.042  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 0.700 4.915 4.180 ;
        RECT  3.115 2.010 4.915 2.410 ;
        RECT  3.080 2.640 3.420 4.180 ;
        RECT  3.115 0.730 3.420 4.180 ;
        RECT  3.080 0.730 3.420 1.070 ;
        RECT  1.640 3.210 3.420 3.490 ;
        RECT  1.640 3.210 1.980 4.105 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.800 -0.400 4.140 1.700 ;
        RECT  2.355 -0.400 2.700 1.040 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.800 2.640 4.140 5.280 ;
        RECT  2.360 3.720 2.700 5.280 ;
        RECT  0.900 3.690 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.110 1.290 1.410 ;
        RECT  0.990 2.070 2.215 2.410 ;
        RECT  0.990 1.110 1.290 2.940 ;
        RECT  0.180 2.640 1.290 2.940 ;
        RECT  0.180 2.640 0.520 4.180 ;
        RECT  1.760 1.240 2.100 1.840 ;
        RECT  1.760 1.540 2.885 1.840 ;
        RECT  2.445 1.540 2.885 1.980 ;
        RECT  2.445 1.540 2.745 2.980 ;
        RECT  1.545 2.640 2.745 2.980 ;
    END
END BUCX4

MACRO BUCX20
    CLASS CORE ;
    FOREIGN BUCX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.743  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.860 0.700 16.255 4.180 ;
        RECT  5.780 1.760 16.255 2.560 ;
        RECT  14.420 0.700 14.760 4.180 ;
        RECT  12.980 0.700 13.320 4.180 ;
        RECT  11.540 0.700 11.880 4.180 ;
        RECT  10.100 0.700 10.440 4.180 ;
        RECT  8.660 0.700 9.000 4.180 ;
        RECT  7.220 0.700 7.560 4.180 ;
        RECT  5.780 0.830 6.120 4.165 ;
        RECT  2.980 3.030 6.120 3.330 ;
        RECT  4.340 3.030 4.680 4.165 ;
        RECT  2.900 3.755 3.240 4.095 ;
        RECT  2.980 3.030 3.240 4.095 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.547  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.800 0.975 2.140 ;
        RECT  0.125 1.640 0.505 2.140 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.140 2.820 15.480 5.280 ;
        RECT  13.690 2.820 14.040 5.280 ;
        RECT  12.260 2.820 12.600 5.280 ;
        RECT  10.820 2.820 11.160 5.280 ;
        RECT  9.380 2.820 9.720 5.280 ;
        RECT  7.930 2.820 8.280 5.280 ;
        RECT  6.500 2.810 6.840 5.280 ;
        RECT  5.060 3.560 5.400 5.280 ;
        RECT  3.620 3.675 3.960 5.280 ;
        RECT  1.690 3.580 2.520 5.280 ;
        RECT  1.690 2.750 2.030 5.280 ;
        RECT  0.190 2.640 0.530 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.140 -0.400 15.480 1.510 ;
        RECT  13.700 -0.400 14.040 1.510 ;
        RECT  12.260 -0.400 12.600 1.510 ;
        RECT  10.820 -0.400 11.160 1.510 ;
        RECT  9.380 -0.400 9.720 1.510 ;
        RECT  7.940 -0.400 8.280 1.510 ;
        RECT  6.500 -0.400 6.840 1.510 ;
        RECT  5.060 -0.400 5.400 1.170 ;
        RECT  3.450 -0.400 3.790 1.165 ;
        RECT  1.690 -0.400 2.030 1.200 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.810 0.700 1.460 1.570 ;
        RECT  1.205 1.930 4.510 2.270 ;
        RECT  1.205 0.700 1.460 4.180 ;
        RECT  0.910 2.640 1.460 4.180 ;
        RECT  2.570 0.865 2.910 1.700 ;
        RECT  4.020 0.790 4.830 1.700 ;
        RECT  2.570 1.400 5.040 1.700 ;
        RECT  4.740 1.400 5.040 2.800 ;
        RECT  2.400 2.500 5.040 2.800 ;
        RECT  2.400 2.500 2.750 2.990 ;
        RECT  1.205 1.930 3.80 2.270 ;
        RECT  2.570 1.400 4.30 1.700 ;
        RECT  2.400 2.500 4.70 2.800 ;
    END
END BUCX20

MACRO BUCX16
    CLASS CORE ;
    FOREIGN BUCX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.397  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.810 2.450 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.755  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  13.340 0.700 13.735 4.180 ;
        RECT  4.700 1.780 13.735 2.480 ;
        RECT  11.900 0.700 12.240 4.180 ;
        RECT  10.460 0.700 10.800 4.180 ;
        RECT  9.020 0.700 9.360 4.180 ;
        RECT  7.580 0.700 7.920 4.180 ;
        RECT  6.140 0.700 6.480 4.180 ;
        RECT  4.700 0.875 5.040 4.180 ;
        RECT  3.260 3.010 5.040 3.310 ;
        RECT  3.260 3.010 3.600 4.165 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 13.860 0.400 ;
        RECT  12.620 -0.400 12.960 1.510 ;
        RECT  11.180 -0.400 11.520 1.510 ;
        RECT  9.740 -0.400 10.080 1.510 ;
        RECT  8.300 -0.400 8.640 1.510 ;
        RECT  6.860 -0.400 7.200 1.510 ;
        RECT  5.420 -0.400 5.760 1.215 ;
        RECT  3.340 -0.400 3.680 1.070 ;
        RECT  1.380 -0.400 1.720 0.950 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 13.860 5.280 ;
        RECT  12.620 2.730 12.960 5.280 ;
        RECT  11.170 2.730 11.520 5.280 ;
        RECT  9.740 2.730 10.080 5.280 ;
        RECT  8.300 2.730 8.640 5.280 ;
        RECT  6.860 2.730 7.200 5.280 ;
        RECT  5.410 2.730 5.760 5.280 ;
        RECT  3.980 3.540 4.320 5.280 ;
        RECT  1.765 3.825 2.880 5.280 ;
        RECT  1.765 2.640 2.105 5.280 ;
        RECT  0.320 2.680 0.660 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.480 1.070 0.820 1.410 ;
        RECT  0.480 1.180 1.380 1.410 ;
        RECT  1.040 1.930 3.995 2.270 ;
        RECT  1.040 1.180 1.380 3.960 ;
        RECT  2.360 0.860 2.700 1.600 ;
        RECT  4.130 0.630 4.470 1.600 ;
        RECT  2.360 1.300 4.470 1.600 ;
        RECT  4.225 0.630 4.470 2.780 ;
        RECT  2.525 2.500 4.470 2.780 ;
        RECT  2.525 2.500 2.865 3.050 ;
        RECT  1.040 1.930 2.30 2.270 ;
        RECT  2.360 1.300 3.70 1.600 ;
    END
END BUCX16

MACRO BUCX12
    CLASS CORE ;
    FOREIGN BUCX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.720  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.960 1.870 10.585 2.470 ;
        RECT  10.190 0.700 10.585 2.470 ;
        RECT  9.470 1.870 9.810 4.180 ;
        RECT  8.750 0.700 9.090 2.470 ;
        RECT  8.030 1.870 8.370 4.180 ;
        RECT  7.310 0.700 7.650 2.470 ;
        RECT  6.640 1.870 6.980 3.450 ;
        RECT  5.870 0.700 6.210 2.470 ;
        RECT  5.300 1.870 5.640 3.450 ;
        RECT  4.430 0.700 4.770 2.470 ;
        RECT  2.570 3.110 4.300 3.450 ;
        RECT  3.960 1.870 4.300 3.450 ;
        RECT  2.570 3.110 2.910 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.101  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.400 0.510 2.210 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.620 ;
        RECT  8.030 -0.400 8.370 1.620 ;
        RECT  6.590 -0.400 6.930 1.620 ;
        RECT  5.150 -0.400 5.490 1.620 ;
        RECT  3.290 -0.400 3.630 1.050 ;
        RECT  1.510 -0.400 1.850 1.220 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 2.740 10.530 5.280 ;
        RECT  8.750 2.725 9.090 5.280 ;
        RECT  7.310 3.640 7.650 5.280 ;
        RECT  5.970 3.640 6.310 5.280 ;
        RECT  4.630 3.640 4.970 5.280 ;
        RECT  3.290 3.680 3.630 5.280 ;
        RECT  0.180 4.160 2.015 5.280 ;
        RECT  1.675 3.220 2.015 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.650 0.790 1.080 1.130 ;
        RECT  0.740 1.830 3.200 2.170 ;
        RECT  0.740 0.790 1.080 3.760 ;
        RECT  2.420 0.790 2.760 1.600 ;
        RECT  3.860 0.730 4.200 1.600 ;
        RECT  2.420 1.300 4.200 1.600 ;
        RECT  3.430 1.300 3.730 2.740 ;
        RECT  2.070 2.400 3.730 2.740 ;
        RECT  0.740 1.830 2.10 2.170 ;
    END
END BUCX12

MACRO BTLX8
    CLASS CORE ;
    FOREIGN BTLX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 5.573  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.815 0.700 11.215 4.180 ;
        RECT  6.490 1.860 11.215 2.360 ;
        RECT  10.810 0.700 11.215 2.360 ;
        RECT  9.375 0.700 9.720 2.360 ;
        RECT  9.375 0.700 9.715 4.180 ;
        RECT  7.935 0.700 8.285 2.360 ;
        RECT  7.935 0.700 8.275 4.180 ;
        RECT  6.490 0.700 6.830 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.716  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.680 4.130 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.458  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.845 2.070 4.660 2.410 ;
        RECT  3.955 2.070 4.285 2.630 ;
        RECT  3.950 2.070 4.285 2.585 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.095 2.640 10.435 5.280 ;
        RECT  8.655 2.590 8.995 5.280 ;
        RECT  7.210 2.590 7.550 5.280 ;
        RECT  5.680 3.355 6.020 5.280 ;
        RECT  4.105 3.320 4.445 5.280 ;
        RECT  1.065 2.740 1.405 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.100 -0.400 10.440 1.575 ;
        RECT  8.660 -0.400 9.000 1.570 ;
        RECT  7.215 -0.400 7.555 1.570 ;
        RECT  5.525 -0.400 5.865 0.940 ;
        RECT  4.045 -0.400 4.385 1.075 ;
        RECT  1.145 -0.400 1.485 1.570 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.170 1.435 2.510 ;
        RECT  0.180 1.175 0.520 3.220 ;
        RECT  1.905 0.630 3.665 0.885 ;
        RECT  3.325 0.630 3.665 1.535 ;
        RECT  3.325 1.305 5.105 1.535 ;
        RECT  4.765 0.700 5.105 1.840 ;
        RECT  4.755 1.305 5.105 1.840 ;
        RECT  4.755 1.585 6.255 1.840 ;
        RECT  5.915 1.170 6.255 1.980 ;
        RECT  1.905 0.630 2.245 2.455 ;
        RECT  1.905 2.225 2.925 2.455 ;
        RECT  2.585 2.225 2.925 3.790 ;
        RECT  2.625 1.150 2.965 1.995 ;
        RECT  2.625 1.765 3.615 1.995 ;
        RECT  3.385 1.765 3.615 4.250 ;
        RECT  3.385 2.860 6.260 3.090 ;
        RECT  5.920 2.310 6.260 3.120 ;
        RECT  4.825 2.590 6.260 3.120 ;
        RECT  1.825 2.685 2.165 4.250 ;
        RECT  4.825 2.590 5.165 4.185 ;
        RECT  3.385 2.635 3.725 4.250 ;
        RECT  1.825 4.020 3.725 4.250 ;
        RECT  3.385 2.860 5.30 3.090 ;
    END
END BTLX8

MACRO BTLX6
    CLASS CORE ;
    FOREIGN BTLX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.122  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.885 0.700 9.325 4.180 ;
        RECT  6.005 1.870 9.325 2.210 ;
        RECT  8.880 0.700 9.325 2.210 ;
        RECT  7.445 0.700 7.790 2.210 ;
        RECT  7.445 0.700 7.785 4.180 ;
        RECT  6.005 0.700 6.355 2.210 ;
        RECT  6.005 0.700 6.345 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.475  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.415 2.595 2.230 2.935 ;
        RECT  1.415 1.610 1.645 2.935 ;
        RECT  0.755 1.610 1.645 2.020 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.895  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.790 1.640 4.285 2.220 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.165 2.740 8.505 5.280 ;
        RECT  6.725 2.740 7.065 5.280 ;
        RECT  5.285 2.730 5.625 5.280 ;
        RECT  3.805 2.945 4.145 5.280 ;
        RECT  0.760 4.050 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.170 -0.400 8.510 1.575 ;
        RECT  6.730 -0.400 7.070 1.570 ;
        RECT  5.285 -0.400 5.625 1.520 ;
        RECT  3.805 -0.400 4.145 1.410 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.280 1.185 2.620 ;
        RECT  0.180 1.090 0.520 3.570 ;
        RECT  1.880 0.630 3.420 0.975 ;
        RECT  1.880 0.630 2.115 1.325 ;
        RECT  1.620 0.985 2.115 1.325 ;
        RECT  3.080 0.630 3.420 1.445 ;
        RECT  1.885 0.630 2.115 2.365 ;
        RECT  1.885 2.135 2.690 2.365 ;
        RECT  2.460 2.135 2.690 3.515 ;
        RECT  2.280 3.170 2.690 3.515 ;
        RECT  2.380 1.360 2.720 1.905 ;
        RECT  2.380 1.675 3.150 1.905 ;
        RECT  2.920 2.485 4.865 2.715 ;
        RECT  2.920 2.485 3.425 3.560 ;
        RECT  4.525 2.485 4.865 3.560 ;
        RECT  1.520 3.195 1.860 4.085 ;
        RECT  2.920 1.675 3.150 4.085 ;
        RECT  1.520 3.745 3.150 4.085 ;
        RECT  4.525 1.105 4.865 2.090 ;
        RECT  4.525 1.750 5.775 2.090 ;
    END
END BTLX6

MACRO BTLX4
    CLASS CORE ;
    FOREIGN BTLX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.945 0.995 7.435 4.120 ;
        RECT  5.505 1.840 7.435 2.530 ;
        RECT  5.505 0.995 5.855 2.530 ;
        RECT  5.505 0.995 5.845 4.120 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.425 2.640 2.050 2.985 ;
        RECT  1.425 1.545 1.655 2.985 ;
        RECT  0.755 1.545 1.655 2.020 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.749  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 1.640 3.885 2.220 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.665 2.800 8.005 5.280 ;
        RECT  6.225 2.800 6.565 5.280 ;
        RECT  4.785 2.800 5.125 5.280 ;
        RECT  3.305 2.910 3.645 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 1.335 ;
        RECT  6.230 -0.400 6.570 1.335 ;
        RECT  4.785 -0.400 5.125 1.335 ;
        RECT  3.305 -0.400 3.645 1.400 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.250 1.195 2.555 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.880 0.785 3.040 1.130 ;
        RECT  1.620 0.975 2.115 1.315 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.615 2.410 ;
        RECT  2.280 2.180 2.615 3.515 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.075 1.950 ;
        RECT  2.845 2.450 4.365 2.680 ;
        RECT  1.520 3.245 1.860 4.085 ;
        RECT  4.025 2.450 4.365 3.865 ;
        RECT  2.845 1.720 3.075 4.085 ;
        RECT  1.520 3.745 3.075 4.085 ;
        RECT  4.025 1.105 4.365 1.450 ;
        RECT  4.115 1.105 4.365 2.110 ;
        RECT  4.115 1.880 5.275 2.110 ;
        RECT  4.935 1.880 5.275 2.220 ;
    END
END BTLX4

MACRO BTLX3
    CLASS CORE ;
    FOREIGN BTLX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.945 0.995 7.435 3.965 ;
        RECT  5.505 1.840 7.435 2.180 ;
        RECT  5.505 0.995 5.855 2.180 ;
        RECT  5.505 0.995 5.845 3.965 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.425 2.640 2.050 2.985 ;
        RECT  1.425 1.545 1.655 2.985 ;
        RECT  0.755 1.545 1.655 2.020 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.567  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 1.635 3.885 2.040 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.225 2.645 6.565 5.280 ;
        RECT  4.785 2.645 5.125 5.280 ;
        RECT  3.305 2.730 3.645 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.230 -0.400 6.570 1.335 ;
        RECT  4.785 -0.400 5.125 1.335 ;
        RECT  3.305 -0.400 3.645 1.400 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.250 1.195 2.555 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  1.880 0.785 3.040 1.130 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.615 2.410 ;
        RECT  2.280 2.180 2.615 3.255 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.075 1.950 ;
        RECT  2.845 2.270 4.365 2.500 ;
        RECT  1.520 3.245 1.860 3.825 ;
        RECT  4.025 2.270 4.365 3.540 ;
        RECT  2.845 1.720 3.075 3.825 ;
        RECT  1.520 3.485 3.075 3.825 ;
        RECT  4.025 1.105 4.365 1.450 ;
        RECT  4.115 1.105 4.365 1.930 ;
        RECT  4.115 1.700 5.275 1.930 ;
        RECT  4.935 1.700 5.275 2.040 ;
    END
END BTLX3

MACRO BTLX20
    CLASS CORE ;
    FOREIGN BTLX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.570 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.493  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  24.050 0.700 24.445 4.180 ;
        RECT  13.925 1.840 24.445 2.490 ;
        RECT  22.610 0.700 22.950 4.180 ;
        RECT  22.600 0.700 22.950 2.490 ;
        RECT  21.170 0.700 21.515 4.180 ;
        RECT  21.160 0.700 21.515 2.490 ;
        RECT  19.730 0.700 20.070 4.180 ;
        RECT  19.725 0.700 20.070 2.490 ;
        RECT  18.290 0.700 18.630 4.180 ;
        RECT  18.285 0.700 18.630 2.490 ;
        RECT  16.850 0.700 17.200 2.490 ;
        RECT  16.850 0.700 17.190 4.180 ;
        RECT  15.405 0.700 15.745 4.180 ;
        RECT  13.965 0.700 14.305 2.490 ;
        RECT  13.925 1.030 14.265 4.180 ;
        RECT  12.445 2.810 14.265 3.110 ;
        RECT  12.445 1.030 14.305 1.330 ;
        RECT  12.445 2.810 12.785 4.180 ;
        RECT  12.445 0.815 12.785 1.330 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.768  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.880 0.530 2.630 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.780  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.750 2.070 7.510 2.410 ;
        RECT  5.845 2.070 6.175 2.630 ;
        RECT  5.830 2.070 6.175 2.590 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 24.570 5.280 ;
        RECT  23.330 2.760 23.670 5.280 ;
        RECT  21.890 2.760 22.230 5.280 ;
        RECT  20.450 2.760 20.790 5.280 ;
        RECT  19.010 2.760 19.350 5.280 ;
        RECT  17.570 2.760 17.910 5.280 ;
        RECT  16.130 2.760 16.470 5.280 ;
        RECT  14.645 2.760 14.985 5.280 ;
        RECT  13.205 3.340 13.545 5.280 ;
        RECT  11.725 2.810 12.065 5.280 ;
        RECT  10.305 2.810 10.645 5.280 ;
        RECT  8.865 2.810 9.205 5.280 ;
        RECT  7.425 3.150 7.765 5.280 ;
        RECT  5.985 3.320 6.325 5.280 ;
        RECT  3.065 3.145 3.405 5.280 ;
        RECT  1.625 2.690 1.965 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 24.570 0.400 ;
        RECT  23.330 -0.400 23.670 1.570 ;
        RECT  21.890 -0.400 22.230 1.570 ;
        RECT  20.450 -0.400 20.790 1.575 ;
        RECT  19.010 -0.400 19.350 1.570 ;
        RECT  17.570 -0.400 17.910 1.570 ;
        RECT  16.125 -0.400 16.465 1.570 ;
        RECT  14.685 -0.400 15.025 1.570 ;
        RECT  13.205 -0.400 13.545 0.800 ;
        RECT  11.725 -0.400 12.065 1.170 ;
        RECT  10.305 -0.400 10.645 1.510 ;
        RECT  8.865 -0.400 9.205 1.510 ;
        RECT  7.425 -0.400 7.765 1.115 ;
        RECT  5.985 -0.400 6.325 1.120 ;
        RECT  3.100 -0.400 3.445 1.315 ;
        RECT  1.625 -0.400 1.970 1.295 ;
        RECT  0.180 -0.400 0.520 1.650 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.120 2.155 2.460 ;
        RECT  0.900 0.830 1.240 3.910 ;
        RECT  4.545 1.115 4.885 1.995 ;
        RECT  4.545 1.765 5.475 1.995 ;
        RECT  8.145 2.240 13.135 2.580 ;
        RECT  5.245 1.765 5.475 4.250 ;
        RECT  2.345 2.685 4.165 2.915 ;
        RECT  6.705 2.690 8.490 2.920 ;
        RECT  5.245 2.860 7.045 3.090 ;
        RECT  2.345 2.685 2.685 3.560 ;
        RECT  3.825 2.685 4.165 4.250 ;
        RECT  6.705 2.690 7.045 4.115 ;
        RECT  8.145 2.240 8.490 4.120 ;
        RECT  9.585 2.240 9.925 4.135 ;
        RECT  11.025 2.240 11.365 4.135 ;
        RECT  5.245 2.640 5.605 4.250 ;
        RECT  3.825 4.020 5.605 4.250 ;
        RECT  3.825 0.630 5.605 0.885 ;
        RECT  5.265 0.630 5.605 1.535 ;
        RECT  6.705 0.740 7.045 1.620 ;
        RECT  5.265 1.305 5.845 1.535 ;
        RECT  2.380 0.975 2.725 1.780 ;
        RECT  11.025 0.940 11.365 1.970 ;
        RECT  5.660 1.390 8.485 1.620 ;
        RECT  8.145 0.740 8.485 1.970 ;
        RECT  8.140 1.390 8.485 1.970 ;
        RECT  9.585 0.740 9.925 1.970 ;
        RECT  2.380 1.550 4.165 1.780 ;
        RECT  11.025 1.560 13.135 1.970 ;
        RECT  8.140 1.740 13.135 1.970 ;
        RECT  3.825 0.630 4.165 2.455 ;
        RECT  3.825 2.225 4.885 2.455 ;
        RECT  4.545 2.225 4.885 3.790 ;
        RECT  8.145 2.240 12.20 2.580 ;
        RECT  5.660 1.390 7.80 1.620 ;
        RECT  11.025 1.560 12.60 1.970 ;
        RECT  8.140 1.740 12.60 1.970 ;
    END
END BTLX20

MACRO BTLX2
    CLASS CORE ;
    FOREIGN BTLX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.425 2.640 2.110 2.985 ;
        RECT  1.425 1.545 1.655 2.985 ;
        RECT  0.755 1.545 1.655 2.020 ;
        END
    END EN
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.192  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.580 1.050 4.920 3.240 ;
        RECT  4.430 2.645 4.770 3.965 ;
        RECT  4.430 1.050 4.920 1.400 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.945 3.655 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 2.645 5.490 5.280 ;
        RECT  3.710 2.860 4.050 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.150 -0.400 5.490 1.070 ;
        RECT  3.705 -0.400 4.045 1.150 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.250 1.195 2.555 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.040 1.950 ;
        RECT  2.810 1.720 3.040 4.105 ;
        RECT  1.520 3.245 1.860 4.105 ;
        RECT  2.810 2.860 3.290 4.105 ;
        RECT  1.520 3.765 3.290 4.105 ;
        RECT  1.880 0.730 3.475 1.070 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  3.245 0.730 3.475 1.610 ;
        RECT  3.245 1.380 4.200 1.610 ;
        RECT  3.970 1.380 4.200 1.970 ;
        RECT  3.970 1.630 4.310 1.970 ;
        RECT  1.885 0.730 2.115 2.410 ;
        RECT  1.885 2.180 2.580 2.410 ;
        RECT  2.350 2.180 2.580 3.525 ;
        RECT  2.240 3.185 2.580 3.525 ;
    END
END BTLX2

MACRO BTLX16
    CLASS CORE ;
    FOREIGN BTLX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 9.557  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.970 0.700 19.405 4.150 ;
        RECT  10.325 1.840 19.405 2.440 ;
        RECT  17.530 0.700 17.870 4.150 ;
        RECT  17.520 0.700 17.870 2.440 ;
        RECT  16.090 0.700 16.435 4.150 ;
        RECT  16.080 0.700 16.435 2.440 ;
        RECT  14.650 0.700 14.990 4.150 ;
        RECT  14.645 0.700 14.990 2.440 ;
        RECT  13.210 0.700 13.550 4.150 ;
        RECT  13.205 0.700 13.550 2.440 ;
        RECT  11.855 1.840 12.195 3.415 ;
        RECT  11.770 0.700 12.120 2.440 ;
        RECT  10.585 1.840 10.925 3.415 ;
        RECT  10.325 0.700 10.665 2.440 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.307  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 1.640 1.200 2.220 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.916  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.025 2.070 6.315 2.410 ;
        RECT  5.165 2.070 5.545 2.630 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.250 -0.400 18.590 1.570 ;
        RECT  16.810 -0.400 17.150 1.570 ;
        RECT  15.370 -0.400 15.710 1.575 ;
        RECT  13.930 -0.400 14.270 1.570 ;
        RECT  12.490 -0.400 12.830 1.570 ;
        RECT  11.045 -0.400 11.385 1.570 ;
        RECT  9.565 -0.400 9.905 1.280 ;
        RECT  8.145 -0.400 8.485 1.510 ;
        RECT  6.705 -0.400 7.045 1.115 ;
        RECT  5.265 -0.400 5.605 1.115 ;
        RECT  2.385 -0.400 2.725 1.410 ;
        RECT  0.905 -0.400 1.245 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.250 2.740 18.590 5.280 ;
        RECT  16.810 2.730 17.150 5.280 ;
        RECT  15.370 2.740 15.710 5.280 ;
        RECT  13.930 2.740 14.270 5.280 ;
        RECT  12.490 3.810 12.830 5.280 ;
        RECT  11.220 3.810 11.560 5.280 ;
        RECT  9.950 3.800 10.290 5.280 ;
        RECT  8.145 2.850 8.485 5.280 ;
        RECT  6.705 3.150 7.045 5.280 ;
        RECT  5.265 3.320 5.605 5.280 ;
        RECT  2.385 3.370 2.725 5.280 ;
        RECT  0.905 2.910 1.245 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.425 2.310 1.765 2.650 ;
        RECT  0.180 2.450 1.545 2.680 ;
        RECT  0.180 0.700 0.520 4.180 ;
        RECT  3.825 1.115 4.165 1.995 ;
        RECT  3.825 1.765 4.775 1.995 ;
        RECT  7.425 2.280 9.000 2.620 ;
        RECT  4.545 1.765 4.775 4.250 ;
        RECT  5.985 2.690 7.765 2.920 ;
        RECT  8.715 2.280 9.000 2.920 ;
        RECT  4.545 2.860 6.325 3.090 ;
        RECT  1.665 2.880 3.445 3.140 ;
        RECT  1.665 2.880 2.005 3.870 ;
        RECT  3.105 2.685 3.445 4.250 ;
        RECT  5.985 2.690 6.325 4.125 ;
        RECT  7.425 2.280 7.765 4.125 ;
        RECT  8.865 2.625 9.715 4.140 ;
        RECT  4.545 2.640 4.885 4.250 ;
        RECT  3.105 4.020 4.885 4.250 ;
        RECT  3.105 0.630 4.885 0.885 ;
        RECT  4.545 0.630 4.885 1.535 ;
        RECT  5.985 0.740 6.325 1.620 ;
        RECT  4.545 1.305 5.135 1.535 ;
        RECT  8.865 0.940 9.210 1.970 ;
        RECT  4.955 1.390 7.765 1.620 ;
        RECT  7.425 0.740 7.765 1.970 ;
        RECT  7.415 1.390 7.765 1.970 ;
        RECT  1.665 1.100 2.005 2.000 ;
        RECT  8.865 1.610 10.045 1.950 ;
        RECT  7.415 1.740 9.570 1.970 ;
        RECT  1.665 1.770 3.445 2.000 ;
        RECT  3.105 0.630 3.445 2.455 ;
        RECT  9.230 1.610 9.570 2.395 ;
        RECT  3.105 2.225 4.165 2.455 ;
        RECT  3.825 2.225 4.165 3.790 ;
        RECT  4.955 1.390 6.90 1.620 ;
        RECT  7.415 1.740 8.80 1.970 ;
    END
END BTLX16

MACRO BTLX12
    CLASS CORE ;
    FOREIGN BTLX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.258  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.140 0.700 15.625 4.180 ;
        RECT  9.375 1.840 15.625 2.390 ;
        RECT  15.130 0.700 15.625 2.390 ;
        RECT  13.700 0.700 14.045 2.390 ;
        RECT  13.700 0.700 14.040 4.180 ;
        RECT  12.260 0.700 12.600 4.180 ;
        RECT  12.255 0.700 12.600 2.390 ;
        RECT  10.820 0.700 11.170 2.390 ;
        RECT  10.820 0.700 11.160 4.180 ;
        RECT  9.375 0.700 9.715 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.091  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 1.640 1.210 2.140 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.272  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.005 2.070 6.295 2.410 ;
        RECT  5.165 2.070 5.545 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.860 2.640 16.200 5.280 ;
        RECT  14.420 2.660 14.760 5.280 ;
        RECT  12.980 2.660 13.320 5.280 ;
        RECT  11.540 2.660 11.880 5.280 ;
        RECT  10.100 2.660 10.440 5.280 ;
        RECT  8.125 2.830 8.955 5.280 ;
        RECT  6.685 3.150 7.025 5.280 ;
        RECT  5.245 3.320 5.585 5.280 ;
        RECT  2.385 3.290 2.725 5.280 ;
        RECT  0.905 2.830 1.245 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.855 -0.400 16.200 1.630 ;
        RECT  14.420 -0.400 14.760 1.575 ;
        RECT  12.980 -0.400 13.320 1.570 ;
        RECT  11.540 -0.400 11.880 1.570 ;
        RECT  10.095 -0.400 10.435 1.570 ;
        RECT  8.165 -0.400 8.505 1.510 ;
        RECT  6.685 -0.400 7.025 1.115 ;
        RECT  5.245 -0.400 5.585 1.115 ;
        RECT  2.385 -0.400 2.725 1.525 ;
        RECT  0.905 -0.400 1.245 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.425 2.230 1.765 2.600 ;
        RECT  0.180 2.370 1.765 2.600 ;
        RECT  0.180 0.810 0.520 3.910 ;
        RECT  3.085 0.795 4.865 1.050 ;
        RECT  4.525 0.795 4.865 1.535 ;
        RECT  5.965 0.740 6.305 1.620 ;
        RECT  4.525 1.305 5.115 1.535 ;
        RECT  4.935 1.390 7.745 1.620 ;
        RECT  7.405 0.740 7.745 1.970 ;
        RECT  7.395 1.390 7.745 1.970 ;
        RECT  1.665 1.215 2.005 2.000 ;
        RECT  8.800 1.140 9.140 1.970 ;
        RECT  7.395 1.740 9.140 1.970 ;
        RECT  1.665 1.770 3.425 2.000 ;
        RECT  3.085 0.795 3.425 2.455 ;
        RECT  3.085 2.225 4.145 2.455 ;
        RECT  3.805 2.225 4.145 3.770 ;
        RECT  3.805 1.280 4.145 1.995 ;
        RECT  3.805 1.765 4.755 1.995 ;
        RECT  7.405 2.280 9.145 2.600 ;
        RECT  4.525 1.765 4.755 4.230 ;
        RECT  5.965 2.690 7.745 2.920 ;
        RECT  1.665 2.830 3.425 3.060 ;
        RECT  4.525 2.860 6.305 3.090 ;
        RECT  1.665 2.830 2.005 3.670 ;
        RECT  3.085 2.830 3.425 4.230 ;
        RECT  5.965 2.690 6.305 4.125 ;
        RECT  7.405 2.280 7.745 4.125 ;
        RECT  4.525 2.640 4.865 4.230 ;
        RECT  3.085 4.000 4.865 4.230 ;
        RECT  4.935 1.390 6.20 1.620 ;
    END
END BTLX12

MACRO BTLX1
    CLASS CORE ;
    FOREIGN BTLX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.425 2.640 2.110 2.985 ;
        RECT  1.425 1.545 1.655 2.985 ;
        RECT  0.755 1.545 1.655 2.020 ;
        END
    END EN
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.056  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.610 0.910 4.925 3.240 ;
        RECT  4.450 2.645 4.790 3.965 ;
        RECT  4.520 0.910 4.925 1.260 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.290 1.640 3.660 2.325 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.720 2.645 4.070 5.280 ;
        RECT  0.780 4.005 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.760 -0.400 4.100 0.710 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.250 1.195 2.555 ;
        RECT  0.180 1.025 0.520 3.505 ;
        RECT  2.380 1.115 2.720 1.950 ;
        RECT  2.380 1.720 3.060 1.950 ;
        RECT  2.830 1.720 3.060 4.075 ;
        RECT  2.830 2.750 3.300 3.090 ;
        RECT  1.540 3.245 1.880 4.075 ;
        RECT  2.830 2.750 3.115 4.075 ;
        RECT  1.540 3.735 3.115 4.075 ;
        RECT  1.880 0.635 3.310 0.865 ;
        RECT  3.080 0.635 3.310 1.410 ;
        RECT  1.880 0.635 2.115 1.315 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  3.080 1.110 4.290 1.410 ;
        RECT  4.040 1.110 4.290 1.970 ;
        RECT  4.040 1.630 4.380 1.970 ;
        RECT  1.885 0.635 2.115 2.410 ;
        RECT  1.885 2.180 2.600 2.410 ;
        RECT  2.370 2.180 2.600 3.505 ;
        RECT  2.260 3.165 2.600 3.505 ;
    END
END BTLX1

MACRO BTLX0
    CLASS CORE ;
    FOREIGN BTLX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.360 2.245 4.285 2.580 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.480 3.320 4.915 3.660 ;
        RECT  4.600 0.910 4.915 3.660 ;
        RECT  4.535 0.910 4.915 1.390 ;
        RECT  4.480 0.910 4.915 1.250 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 2.105 2.200 2.795 ;
        RECT  1.860 2.105 2.195 2.800 ;
        RECT  0.755 2.105 2.200 2.335 ;
        RECT  0.755 1.535 1.135 2.335 ;
        END
    END EN
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.680 4.060 4.020 5.280 ;
        RECT  0.780 3.770 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.815 -0.400 4.120 0.710 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.565 1.470 2.845 ;
        RECT  0.180 1.110 0.520 3.370 ;
        RECT  2.380 1.165 3.125 1.415 ;
        RECT  2.895 1.165 3.125 3.040 ;
        RECT  3.080 2.810 4.370 3.095 ;
        RECT  1.580 3.050 1.920 3.730 ;
        RECT  3.080 2.810 3.420 3.730 ;
        RECT  1.580 3.500 3.420 3.730 ;
        RECT  1.580 0.650 3.585 0.935 ;
        RECT  3.355 0.650 3.585 1.875 ;
        RECT  1.580 0.650 1.920 1.875 ;
        RECT  1.580 1.645 2.665 1.875 ;
        RECT  3.355 1.560 4.370 1.875 ;
        RECT  2.435 1.645 2.665 3.270 ;
        RECT  2.385 2.935 2.665 3.270 ;
        RECT  1.580 0.650 2.80 0.935 ;
    END
END BTLX0

MACRO BTLCX8
    CLASS CORE ;
    FOREIGN BTLCX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 5.101  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.835 1.925 10.585 2.265 ;
        RECT  10.190 0.700 10.585 2.265 ;
        RECT  7.310 1.765 10.585 2.265 ;
        RECT  9.470 1.765 9.810 4.180 ;
        RECT  8.750 0.700 9.090 2.265 ;
        RECT  8.030 1.765 8.370 3.430 ;
        RECT  7.310 0.700 7.650 2.265 ;
        RECT  5.870 1.270 7.650 1.500 ;
        RECT  6.690 2.620 7.115 3.430 ;
        RECT  6.835 1.925 7.115 3.430 ;
        RECT  5.350 2.830 7.115 3.170 ;
        RECT  5.870 0.700 6.210 1.500 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.747  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.920 1.640 3.260 1.980 ;
        RECT  0.655 1.640 3.260 1.890 ;
        RECT  0.655 1.640 1.135 2.020 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.934  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.880 1.640 5.545 2.100 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 2.640 10.530 5.280 ;
        RECT  8.750 2.620 9.090 5.280 ;
        RECT  7.360 3.620 7.700 5.280 ;
        RECT  6.020 3.660 6.360 5.280 ;
        RECT  3.580 3.910 3.920 5.280 ;
        RECT  2.060 3.960 2.400 5.280 ;
        RECT  0.940 3.960 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.535 ;
        RECT  8.030 -0.400 8.370 1.535 ;
        RECT  6.590 -0.400 6.930 1.040 ;
        RECT  5.150 -0.400 5.490 1.275 ;
        RECT  3.430 -0.400 3.770 0.710 ;
        RECT  1.480 -0.400 1.820 1.365 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.170 0.905 1.060 1.245 ;
        RECT  0.170 0.905 0.400 3.560 ;
        RECT  1.790 2.120 2.130 2.480 ;
        RECT  0.170 2.250 2.130 2.480 ;
        RECT  0.170 2.250 0.520 3.560 ;
        RECT  2.730 0.955 4.080 1.295 ;
        RECT  1.500 2.710 4.080 3.005 ;
        RECT  3.780 0.955 4.080 3.680 ;
        RECT  1.500 2.710 1.840 3.560 ;
        RECT  2.820 2.710 3.160 3.560 ;
        RECT  3.780 3.400 5.280 3.680 ;
        RECT  4.940 3.400 5.280 4.250 ;
        RECT  5.795 1.730 6.605 2.070 ;
        RECT  4.310 0.700 4.650 2.600 ;
        RECT  5.795 1.730 6.065 2.600 ;
        RECT  4.310 2.330 6.065 2.600 ;
        RECT  4.570 2.330 4.910 3.170 ;
        RECT  1.500 2.710 3.30 3.005 ;
    END
END BTLCX8

MACRO BTLCX6
    CLASS CORE ;
    FOREIGN BTLCX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.035  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.985 1.830 8.695 2.170 ;
        RECT  8.145 1.640 8.695 2.170 ;
        RECT  8.145 0.700 8.485 2.170 ;
        RECT  7.425 1.830 7.765 4.190 ;
        RECT  6.705 0.700 7.045 2.170 ;
        RECT  5.985 1.310 6.325 4.170 ;
        RECT  4.545 2.790 6.325 3.090 ;
        RECT  5.265 1.310 6.325 1.610 ;
        RECT  5.265 0.700 5.605 1.610 ;
        RECT  4.545 2.790 4.885 4.170 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.614  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.590 1.625 2.580 1.965 ;
        RECT  0.590 1.625 1.135 2.020 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.877  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.155 1.640 4.890 2.030 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.145 2.640 8.485 5.280 ;
        RECT  6.705 2.640 7.045 5.280 ;
        RECT  5.265 3.320 5.605 5.280 ;
        RECT  3.710 3.830 4.050 5.280 ;
        RECT  2.220 2.740 2.565 5.280 ;
        RECT  0.780 3.460 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.425 -0.400 7.765 1.580 ;
        RECT  5.985 -0.400 6.325 1.080 ;
        RECT  4.545 -0.400 4.885 1.275 ;
        RECT  2.765 -0.400 3.105 0.710 ;
        RECT  0.780 -0.400 1.120 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.130 1.025 0.520 1.365 ;
        RECT  0.130 1.025 0.360 4.250 ;
        RECT  0.130 2.680 0.520 4.250 ;
        RECT  2.050 0.985 3.140 1.325 ;
        RECT  1.500 2.210 3.140 2.510 ;
        RECT  2.840 0.985 3.140 3.600 ;
        RECT  2.840 3.260 4.290 3.600 ;
        RECT  1.500 2.210 1.840 4.180 ;
        RECT  3.430 0.935 4.025 1.275 ;
        RECT  3.430 0.935 3.775 2.560 ;
        RECT  5.120 1.840 5.460 2.560 ;
        RECT  3.430 2.260 5.460 2.560 ;
        RECT  3.430 0.935 3.770 3.030 ;
        RECT  3.430 2.260 4.70 2.560 ;
    END
END BTLCX6

MACRO BTLCX4
    CLASS CORE ;
    FOREIGN BTLCX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.649  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 1.640 6.750 2.040 ;
        RECT  6.410 0.700 6.750 2.040 ;
        RECT  5.690 1.640 6.030 4.190 ;
        RECT  4.510 3.240 6.030 3.580 ;
        RECT  5.145 1.010 5.445 2.040 ;
        RECT  4.970 1.010 5.445 1.350 ;
        RECT  4.250 3.740 4.740 4.080 ;
        RECT  4.510 3.240 4.740 4.080 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.437  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.630 1.625 2.580 1.965 ;
        RECT  0.630 1.625 1.135 2.020 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.690  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.440 1.640 4.915 2.020 ;
        RECT  4.440 0.940 4.740 2.020 ;
        RECT  3.650 0.940 4.740 1.170 ;
        RECT  3.650 0.645 3.980 1.170 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 2.640 6.750 5.280 ;
        RECT  4.970 3.840 5.310 5.280 ;
        RECT  3.530 3.740 3.870 5.280 ;
        RECT  2.220 2.725 2.565 5.280 ;
        RECT  0.780 3.460 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.370 ;
        RECT  4.210 -0.400 4.550 0.710 ;
        RECT  2.765 -0.400 3.105 0.710 ;
        RECT  0.780 -0.400 1.120 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.170 1.025 0.520 1.365 ;
        RECT  0.170 1.025 0.400 4.250 ;
        RECT  0.170 2.680 0.520 4.250 ;
        RECT  3.410 1.400 3.780 2.685 ;
        RECT  3.410 2.345 4.275 2.685 ;
        RECT  3.410 1.400 3.710 2.980 ;
        RECT  2.050 0.985 3.140 1.325 ;
        RECT  1.500 2.195 3.140 2.495 ;
        RECT  2.840 0.985 3.140 3.510 ;
        RECT  3.940 3.015 4.280 3.510 ;
        RECT  2.840 3.210 4.280 3.510 ;
        RECT  1.500 2.195 1.840 4.180 ;
    END
END BTLCX4

MACRO BTLCX20
    CLASS CORE ;
    FOREIGN BTLCX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 11.831  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.380 1.810 18.720 4.130 ;
        RECT  8.945 1.810 18.720 2.460 ;
        RECT  17.650 0.700 18.145 2.460 ;
        RECT  17.000 1.810 17.340 3.370 ;
        RECT  16.210 0.700 16.550 2.460 ;
        RECT  15.720 1.810 16.060 3.370 ;
        RECT  14.770 0.700 15.110 2.460 ;
        RECT  14.440 1.810 14.780 3.365 ;
        RECT  13.330 0.700 13.670 2.460 ;
        RECT  13.160 1.810 13.500 3.370 ;
        RECT  11.890 0.700 12.230 2.460 ;
        RECT  11.800 1.810 12.140 4.180 ;
        RECT  10.450 0.700 10.790 2.460 ;
        RECT  10.360 1.810 10.700 4.180 ;
        RECT  8.945 1.340 9.350 2.460 ;
        RECT  9.010 0.700 9.350 2.460 ;
        RECT  8.920 2.390 9.260 4.180 ;
        RECT  7.570 1.340 9.350 1.570 ;
        RECT  7.480 2.390 9.260 2.645 ;
        RECT  7.570 0.700 7.910 1.570 ;
        RECT  7.480 2.390 7.820 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.276  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.440 1.690 3.780 2.030 ;
        RECT  0.755 1.690 3.780 1.920 ;
        RECT  0.755 1.690 1.320 2.220 ;
        RECT  0.755 1.640 1.135 2.220 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.531  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.395 5.585 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  17.660 3.580 18.000 5.280 ;
        RECT  16.360 3.630 16.700 5.280 ;
        RECT  15.080 3.600 15.420 5.280 ;
        RECT  13.800 3.590 14.140 5.280 ;
        RECT  12.520 3.590 12.860 5.280 ;
        RECT  11.080 2.690 11.420 5.280 ;
        RECT  9.640 2.690 9.980 5.280 ;
        RECT  8.200 2.875 8.540 5.280 ;
        RECT  6.760 2.690 7.100 5.280 ;
        RECT  4.220 3.245 4.560 5.280 ;
        RECT  2.780 3.200 3.120 5.280 ;
        RECT  0.180 3.960 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  18.375 -0.400 18.715 1.580 ;
        RECT  16.930 -0.400 17.270 1.580 ;
        RECT  15.490 -0.400 15.830 1.580 ;
        RECT  14.050 -0.400 14.390 1.580 ;
        RECT  12.610 -0.400 12.950 1.580 ;
        RECT  11.170 -0.400 11.510 1.580 ;
        RECT  9.730 -0.400 10.070 1.580 ;
        RECT  8.290 -0.400 8.630 1.110 ;
        RECT  6.850 -0.400 7.190 1.320 ;
        RECT  5.110 -0.400 5.450 1.165 ;
        RECT  3.330 -0.400 3.670 0.710 ;
        RECT  1.500 -0.400 1.840 1.460 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.225 1.120 1.080 1.410 ;
        RECT  0.225 1.120 0.525 2.750 ;
        RECT  1.590 2.150 2.150 2.460 ;
        RECT  0.225 2.450 1.830 2.750 ;
        RECT  0.740 2.450 1.080 3.560 ;
        RECT  2.790 1.075 3.130 1.460 ;
        RECT  2.790 1.230 4.310 1.460 ;
        RECT  4.010 1.230 4.310 3.015 ;
        RECT  2.060 2.690 4.310 2.970 ;
        RECT  3.500 2.785 5.180 3.015 ;
        RECT  4.880 2.785 5.180 4.250 ;
        RECT  6.225 2.700 6.530 4.250 ;
        RECT  2.060 2.690 2.400 4.180 ;
        RECT  3.500 2.690 3.850 4.180 ;
        RECT  6.280 2.500 6.530 4.250 ;
        RECT  4.880 3.950 6.530 4.250 ;
        RECT  4.240 0.700 4.860 1.000 ;
        RECT  5.980 0.825 6.320 2.140 ;
        RECT  5.815 1.800 8.715 2.140 ;
        RECT  4.560 0.700 4.860 2.550 ;
        RECT  5.815 1.800 6.045 2.550 ;
        RECT  4.560 2.250 6.045 2.550 ;
        RECT  5.410 2.250 5.750 3.720 ;
        RECT  2.060 2.690 3.30 2.970 ;
        RECT  5.815 1.800 7.70 2.140 ;
    END
END BTLCX20

MACRO BTLCX16
    CLASS CORE ;
    FOREIGN BTLCX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 10.360  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 0.700 16.885 4.180 ;
        RECT  9.290 1.830 16.885 2.430 ;
        RECT  15.050 0.700 15.390 4.180 ;
        RECT  13.610 0.700 13.950 4.180 ;
        RECT  12.170 0.700 12.510 4.180 ;
        RECT  10.730 0.700 11.070 4.180 ;
        RECT  9.290 0.700 9.630 4.180 ;
        RECT  7.850 2.350 9.630 2.600 ;
        RECT  7.850 1.320 9.630 1.550 ;
        RECT  7.850 2.350 8.190 4.180 ;
        RECT  7.850 0.700 8.190 1.550 ;
        RECT  6.460 2.780 8.190 3.120 ;
        RECT  6.460 2.780 6.750 4.180 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.242  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.320 1.640 3.660 2.030 ;
        RECT  0.755 1.640 3.660 1.890 ;
        RECT  0.755 1.640 1.300 2.030 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.414  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.470 6.070 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 2.660 16.110 5.280 ;
        RECT  14.330 2.660 14.670 5.280 ;
        RECT  12.890 2.660 13.230 5.280 ;
        RECT  11.450 2.660 11.790 5.280 ;
        RECT  10.010 2.660 10.350 5.280 ;
        RECT  8.570 2.830 8.910 5.280 ;
        RECT  7.130 3.350 7.470 5.280 ;
        RECT  4.140 3.245 4.480 5.280 ;
        RECT  2.620 4.170 2.960 5.280 ;
        RECT  0.180 3.830 1.680 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.770 -0.400 16.110 1.600 ;
        RECT  14.330 -0.400 14.670 1.600 ;
        RECT  12.890 -0.400 13.230 1.600 ;
        RECT  11.450 -0.400 11.790 1.600 ;
        RECT  10.010 -0.400 10.350 1.600 ;
        RECT  8.570 -0.400 8.910 1.090 ;
        RECT  7.130 -0.400 7.470 1.165 ;
        RECT  5.250 -0.400 5.590 1.165 ;
        RECT  3.330 -0.400 3.670 0.710 ;
        RECT  1.560 -0.400 1.900 1.320 ;
        RECT  0.240 -0.400 0.580 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.225 1.070 1.180 1.410 ;
        RECT  0.225 1.070 0.525 2.560 ;
        RECT  1.635 2.120 2.160 2.460 ;
        RECT  0.225 2.260 1.865 2.560 ;
        RECT  0.740 2.260 1.080 3.195 ;
        RECT  2.790 1.070 3.130 1.410 ;
        RECT  2.790 1.180 4.120 1.410 ;
        RECT  3.890 1.180 4.120 3.015 ;
        RECT  2.060 2.690 4.120 2.985 ;
        RECT  3.420 2.785 5.010 3.015 ;
        RECT  2.060 2.690 2.400 3.740 ;
        RECT  4.710 2.785 5.010 4.250 ;
        RECT  3.420 2.690 3.770 4.180 ;
        RECT  5.890 2.970 6.230 4.250 ;
        RECT  4.710 3.910 6.230 4.250 ;
        RECT  4.310 0.700 4.650 1.040 ;
        RECT  6.190 0.825 6.600 1.165 ;
        RECT  6.300 1.780 8.890 2.120 ;
        RECT  4.350 0.700 4.650 2.550 ;
        RECT  6.300 0.825 6.600 2.550 ;
        RECT  4.350 2.250 6.600 2.550 ;
        RECT  5.330 2.250 5.660 3.660 ;
        RECT  2.060 2.690 3.90 2.985 ;
        RECT  6.300 1.780 7.70 2.120 ;
        RECT  4.350 2.250 5.80 2.550 ;
    END
END BTLCX16

MACRO BTLCX12
    CLASS CORE ;
    FOREIGN BTLCX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.416  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 1.640 12.475 4.180 ;
        RECT  6.675 1.830 12.475 2.380 ;
        RECT  11.360 1.640 12.475 2.380 ;
        RECT  11.360 0.700 11.700 2.380 ;
        RECT  10.690 1.830 11.030 3.430 ;
        RECT  9.920 0.700 10.260 2.380 ;
        RECT  9.350 1.830 9.690 3.430 ;
        RECT  8.480 0.700 8.820 2.380 ;
        RECT  8.010 1.830 8.350 3.430 ;
        RECT  6.675 1.270 7.380 2.380 ;
        RECT  7.040 0.700 7.380 2.380 ;
        RECT  6.675 1.270 7.015 3.430 ;
        RECT  5.290 2.910 7.015 3.210 ;
        RECT  5.600 1.270 7.380 1.535 ;
        RECT  5.600 0.700 5.940 1.535 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.931  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.780 1.640 3.120 1.985 ;
        RECT  0.755 1.640 3.120 1.890 ;
        RECT  0.755 1.640 1.180 2.030 ;
        END
    END EN
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.020 2.220 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.360 3.620 11.700 5.280 ;
        RECT  10.020 3.620 10.360 5.280 ;
        RECT  8.680 3.620 9.020 5.280 ;
        RECT  7.340 3.625 7.680 5.280 ;
        RECT  6.010 3.660 6.350 5.280 ;
        RECT  3.580 3.910 3.920 5.280 ;
        RECT  2.060 4.170 2.400 5.280 ;
        RECT  0.940 4.170 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.080 -0.400 12.420 1.310 ;
        RECT  10.640 -0.400 10.980 1.580 ;
        RECT  9.200 -0.400 9.540 1.580 ;
        RECT  7.760 -0.400 8.100 1.580 ;
        RECT  6.320 -0.400 6.660 1.040 ;
        RECT  4.880 -0.400 5.220 1.310 ;
        RECT  3.100 -0.400 3.440 0.710 ;
        RECT  1.360 -0.400 1.700 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.905 0.940 1.245 ;
        RECT  1.660 2.120 2.000 2.490 ;
        RECT  0.180 2.260 2.000 2.490 ;
        RECT  0.180 0.905 0.520 3.910 ;
        RECT  2.590 1.070 3.655 1.410 ;
        RECT  3.355 1.070 3.655 3.015 ;
        RECT  1.500 2.720 3.655 3.015 ;
        RECT  2.820 2.720 3.160 3.680 ;
        RECT  2.820 3.440 5.270 3.680 ;
        RECT  1.500 2.720 1.840 3.760 ;
        RECT  4.930 3.440 5.270 4.250 ;
        RECT  4.010 0.700 4.345 1.510 ;
        RECT  5.315 1.765 6.125 2.105 ;
        RECT  4.010 0.700 4.305 2.680 ;
        RECT  5.315 1.765 5.655 2.680 ;
        RECT  4.010 2.450 5.655 2.680 ;
        RECT  4.570 2.450 4.910 3.210 ;
        RECT  1.500 2.720 2.30 3.015 ;
        RECT  2.820 3.440 4.20 3.680 ;
    END
END BTLCX12

MACRO BTHX8
    CLASS CORE ;
    FOREIGN BTHX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.458  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.685 2.070 4.500 2.410 ;
        RECT  3.905 2.070 4.285 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 5.573  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  10.815 0.700 11.215 4.180 ;
        RECT  6.490 1.910 11.215 2.410 ;
        RECT  10.810 0.700 11.215 2.410 ;
        RECT  9.375 0.700 9.720 2.410 ;
        RECT  9.375 0.700 9.715 4.180 ;
        RECT  7.935 0.700 8.285 2.410 ;
        RECT  7.935 0.700 8.275 4.180 ;
        RECT  6.490 0.700 6.830 4.180 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.761  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.680 4.080 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 11.340 0.400 ;
        RECT  10.100 -0.400 10.440 1.635 ;
        RECT  8.660 -0.400 9.000 1.630 ;
        RECT  7.215 -0.400 7.555 1.630 ;
        RECT  5.325 -0.400 5.665 1.330 ;
        RECT  3.885 -0.400 4.225 1.075 ;
        RECT  1.025 -0.400 1.365 1.570 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 11.340 5.280 ;
        RECT  10.095 2.640 10.435 5.280 ;
        RECT  8.655 2.640 8.995 5.280 ;
        RECT  7.210 2.640 7.550 5.280 ;
        RECT  5.385 3.570 6.070 5.280 ;
        RECT  5.385 3.100 5.690 5.280 ;
        RECT  3.945 3.320 4.285 5.280 ;
        RECT  0.945 2.690 1.285 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.800 1.435 2.140 ;
        RECT  0.180 1.175 0.520 3.220 ;
        RECT  1.745 0.630 3.505 0.885 ;
        RECT  3.165 0.630 3.505 1.535 ;
        RECT  3.165 1.305 4.945 1.535 ;
        RECT  4.605 0.700 4.945 1.840 ;
        RECT  4.595 1.305 4.945 1.840 ;
        RECT  4.595 1.560 6.255 1.840 ;
        RECT  5.915 1.170 6.255 1.980 ;
        RECT  1.745 0.630 2.085 2.455 ;
        RECT  1.745 2.225 2.765 2.455 ;
        RECT  2.425 2.225 2.765 3.790 ;
        RECT  2.465 1.150 2.805 1.995 ;
        RECT  2.465 1.765 3.455 1.995 ;
        RECT  3.225 1.765 3.455 4.250 ;
        RECT  4.665 2.590 6.260 2.870 ;
        RECT  3.225 2.860 5.005 3.090 ;
        RECT  5.920 2.310 6.260 3.120 ;
        RECT  1.665 2.685 2.005 4.250 ;
        RECT  4.665 2.590 5.005 4.185 ;
        RECT  3.225 2.635 3.565 4.250 ;
        RECT  1.665 4.020 3.565 4.250 ;
    END
END BTHX8

MACRO BTHX6
    CLASS CORE ;
    FOREIGN BTHX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.895  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.820 1.640 4.340 2.220 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.122  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.930 0.700 9.325 4.180 ;
        RECT  6.050 2.010 9.325 2.350 ;
        RECT  8.920 0.700 9.325 2.350 ;
        RECT  7.490 0.700 7.830 4.180 ;
        RECT  7.485 0.700 7.830 2.350 ;
        RECT  6.050 0.700 6.400 2.350 ;
        RECT  6.050 0.700 6.390 4.180 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.513  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.180 1.135 2.820 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.210 2.640 8.550 5.280 ;
        RECT  6.770 2.640 7.110 5.280 ;
        RECT  5.330 2.640 5.670 5.280 ;
        RECT  3.850 2.945 4.190 5.280 ;
        RECT  0.800 3.720 1.150 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.210 -0.400 8.550 1.575 ;
        RECT  6.770 -0.400 7.110 1.570 ;
        RECT  5.330 -0.400 5.670 1.520 ;
        RECT  3.850 -0.400 4.190 1.410 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.610 1.595 1.950 ;
        RECT  1.365 1.610 1.595 2.940 ;
        RECT  1.365 2.595 2.230 2.940 ;
        RECT  0.180 1.090 0.520 3.280 ;
        RECT  1.880 0.630 3.465 0.975 ;
        RECT  1.620 0.900 2.115 1.240 ;
        RECT  3.125 0.630 3.465 1.445 ;
        RECT  1.885 0.630 2.115 2.365 ;
        RECT  1.885 2.135 2.690 2.365 ;
        RECT  2.460 2.135 2.690 3.515 ;
        RECT  2.280 3.170 2.690 3.515 ;
        RECT  2.380 1.360 2.720 1.905 ;
        RECT  2.380 1.675 3.360 1.905 ;
        RECT  3.130 1.675 3.360 4.085 ;
        RECT  3.130 2.485 4.910 2.715 ;
        RECT  4.570 2.485 4.910 3.560 ;
        RECT  1.520 3.170 1.860 4.085 ;
        RECT  3.130 2.485 3.470 4.085 ;
        RECT  1.520 3.745 3.470 4.085 ;
        RECT  4.570 1.105 4.910 2.090 ;
        RECT  4.570 1.750 5.820 2.090 ;
    END
END BTHX6

MACRO BTHX4
    CLASS CORE ;
    FOREIGN BTHX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.749  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 1.640 3.885 2.220 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.945 0.995 7.435 4.120 ;
        RECT  5.505 2.130 7.435 2.470 ;
        RECT  5.505 0.995 5.855 2.470 ;
        RECT  5.505 0.995 5.845 4.120 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.135 2.890 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.665 2.800 8.005 5.280 ;
        RECT  6.225 2.800 6.565 5.280 ;
        RECT  4.785 2.800 5.125 5.280 ;
        RECT  3.305 2.910 3.645 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.670 -0.400 8.010 1.335 ;
        RECT  6.230 -0.400 6.570 1.335 ;
        RECT  4.785 -0.400 5.125 1.335 ;
        RECT  3.305 -0.400 3.645 1.400 ;
        RECT  0.860 -0.400 1.200 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.050 2.985 ;
        RECT  0.180 1.025 0.520 3.545 ;
        RECT  1.620 0.785 3.040 1.130 ;
        RECT  1.620 0.785 2.115 1.245 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.615 2.410 ;
        RECT  2.280 2.180 2.615 3.515 ;
        RECT  2.380 1.360 3.075 1.700 ;
        RECT  2.845 2.450 4.365 2.680 ;
        RECT  1.520 3.215 1.860 4.085 ;
        RECT  4.025 2.450 4.365 3.865 ;
        RECT  2.845 1.360 3.075 4.085 ;
        RECT  1.520 3.745 3.075 4.085 ;
        RECT  4.025 1.105 4.365 1.450 ;
        RECT  4.115 1.105 4.365 2.110 ;
        RECT  4.115 1.880 5.275 2.110 ;
        RECT  4.935 1.880 5.275 2.220 ;
    END
END BTHX4

MACRO BTHX3
    CLASS CORE ;
    FOREIGN BTHX3 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.567  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.305 1.635 3.885 2.040 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 0.990 7.435 3.965 ;
        RECT  5.600 1.965 7.435 2.305 ;
        RECT  7.035 0.990 7.435 2.305 ;
        RECT  5.600 0.990 5.940 3.965 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.115 1.135 2.755 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 2.645 6.660 5.280 ;
        RECT  4.875 2.645 5.215 5.280 ;
        RECT  3.395 2.730 3.735 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.330 ;
        RECT  4.875 -0.400 5.215 1.330 ;
        RECT  3.395 -0.400 3.735 1.405 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.050 2.985 ;
        RECT  0.180 1.025 0.520 3.545 ;
        RECT  1.880 0.785 3.040 1.130 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  1.885 0.785 2.115 2.410 ;
        RECT  1.885 2.180 2.615 2.410 ;
        RECT  2.280 2.180 2.615 3.255 ;
        RECT  2.380 1.360 3.075 1.700 ;
        RECT  2.845 2.270 4.455 2.500 ;
        RECT  1.520 3.245 1.860 3.825 ;
        RECT  4.115 2.270 4.455 3.540 ;
        RECT  2.845 1.360 3.075 3.825 ;
        RECT  1.520 3.485 3.075 3.825 ;
        RECT  4.115 1.060 4.455 2.040 ;
        RECT  4.115 1.700 5.370 2.040 ;
    END
END BTHX3

MACRO BTHX20
    CLASS CORE ;
    FOREIGN BTHX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.570 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 3.780  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.750 2.070 7.510 2.410 ;
        RECT  5.815 2.070 6.175 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.493  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  24.050 0.700 24.445 4.180 ;
        RECT  13.925 1.840 24.445 2.490 ;
        RECT  22.610 0.700 22.950 4.180 ;
        RECT  22.600 0.700 22.950 2.490 ;
        RECT  21.170 0.700 21.515 4.180 ;
        RECT  21.160 0.700 21.515 2.490 ;
        RECT  19.730 0.700 20.070 4.180 ;
        RECT  19.725 0.700 20.070 2.490 ;
        RECT  18.290 0.700 18.630 4.180 ;
        RECT  18.285 0.700 18.630 2.490 ;
        RECT  16.850 0.700 17.200 2.490 ;
        RECT  16.850 0.700 17.190 4.180 ;
        RECT  15.405 0.700 15.745 4.180 ;
        RECT  13.965 0.700 14.305 2.490 ;
        RECT  13.925 1.030 14.265 4.180 ;
        RECT  12.445 2.810 14.265 3.110 ;
        RECT  12.445 1.030 14.305 1.330 ;
        RECT  12.445 2.810 12.785 4.180 ;
        RECT  12.445 0.815 12.785 1.330 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.721  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.880 0.530 2.630 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 24.570 0.400 ;
        RECT  23.330 -0.400 23.670 1.570 ;
        RECT  21.890 -0.400 22.230 1.570 ;
        RECT  20.450 -0.400 20.790 1.575 ;
        RECT  19.010 -0.400 19.350 1.570 ;
        RECT  17.570 -0.400 17.910 1.570 ;
        RECT  16.125 -0.400 16.465 1.570 ;
        RECT  14.685 -0.400 15.025 1.570 ;
        RECT  13.205 -0.400 13.545 0.800 ;
        RECT  11.725 -0.400 12.065 1.170 ;
        RECT  10.305 -0.400 10.645 1.510 ;
        RECT  8.865 -0.400 9.205 1.510 ;
        RECT  7.425 -0.400 7.765 1.115 ;
        RECT  5.985 -0.400 6.325 1.120 ;
        RECT  3.105 -0.400 3.445 1.555 ;
        RECT  1.625 -0.400 1.965 1.560 ;
        RECT  0.180 -0.400 0.520 1.650 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 24.570 5.280 ;
        RECT  23.330 2.760 23.670 5.280 ;
        RECT  21.890 2.760 22.230 5.280 ;
        RECT  20.450 2.760 20.790 5.280 ;
        RECT  19.010 2.760 19.350 5.280 ;
        RECT  17.570 2.760 17.910 5.280 ;
        RECT  16.130 2.760 16.470 5.280 ;
        RECT  14.645 2.760 14.985 5.280 ;
        RECT  13.205 3.340 13.545 5.280 ;
        RECT  11.725 2.810 12.065 5.280 ;
        RECT  10.305 2.810 10.645 5.280 ;
        RECT  8.865 2.810 9.205 5.280 ;
        RECT  7.425 3.150 7.765 5.280 ;
        RECT  5.985 3.320 6.325 5.280 ;
        RECT  3.105 3.145 3.445 5.280 ;
        RECT  1.625 2.690 2.005 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 1.870 2.155 2.210 ;
        RECT  0.900 0.830 1.240 3.910 ;
        RECT  4.545 1.115 4.885 1.995 ;
        RECT  4.545 1.765 5.475 1.995 ;
        RECT  8.145 2.240 13.135 2.580 ;
        RECT  5.245 1.765 5.475 4.250 ;
        RECT  2.385 2.685 4.145 2.915 ;
        RECT  6.705 2.690 8.490 2.920 ;
        RECT  5.245 2.860 7.045 3.090 ;
        RECT  3.805 2.685 4.145 4.250 ;
        RECT  6.705 2.690 7.045 4.115 ;
        RECT  8.145 2.240 8.490 4.120 ;
        RECT  9.585 2.240 9.925 4.135 ;
        RECT  11.025 2.240 11.365 4.135 ;
        RECT  2.385 2.685 2.725 4.180 ;
        RECT  5.245 2.640 5.585 4.250 ;
        RECT  3.805 4.020 5.585 4.250 ;
        RECT  3.825 0.630 5.605 0.885 ;
        RECT  5.265 0.630 5.605 1.535 ;
        RECT  6.705 0.740 7.045 1.620 ;
        RECT  5.265 1.305 5.845 1.535 ;
        RECT  11.025 0.940 11.365 1.970 ;
        RECT  5.660 1.390 8.485 1.620 ;
        RECT  8.145 0.740 8.485 1.970 ;
        RECT  8.140 1.390 8.485 1.970 ;
        RECT  9.585 0.740 9.925 1.970 ;
        RECT  11.025 1.560 13.135 1.970 ;
        RECT  8.140 1.740 13.135 1.970 ;
        RECT  2.385 1.215 2.725 2.455 ;
        RECT  3.825 0.630 4.165 2.455 ;
        RECT  2.385 2.225 4.865 2.455 ;
        RECT  4.525 2.225 4.865 3.790 ;
        RECT  8.145 2.240 12.80 2.580 ;
        RECT  5.660 1.390 7.60 1.620 ;
        RECT  11.025 1.560 12.40 1.970 ;
        RECT  8.140 1.740 12.90 1.970 ;
        RECT  2.385 2.225 3.40 2.455 ;
    END
END BTHX20

MACRO BTHX2
    CLASS CORE ;
    FOREIGN BTHX2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.945 3.655 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.192  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.580 0.920 4.920 3.240 ;
        RECT  4.430 2.645 4.770 3.965 ;
        RECT  4.430 0.920 4.920 1.270 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.115 1.135 2.755 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 2.645 5.490 5.280 ;
        RECT  3.710 2.860 4.050 5.280 ;
        RECT  0.760 4.005 1.110 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.150 -0.400 5.490 1.260 ;
        RECT  3.705 -0.400 4.045 1.150 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.090 2.985 ;
        RECT  0.180 1.025 0.520 3.545 ;
        RECT  2.380 1.360 2.720 1.950 ;
        RECT  2.380 1.720 3.040 1.950 ;
        RECT  2.810 1.720 3.040 4.105 ;
        RECT  1.520 3.245 1.860 4.105 ;
        RECT  2.810 2.860 3.290 4.105 ;
        RECT  1.520 3.765 3.290 4.105 ;
        RECT  1.880 0.730 3.475 1.070 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  3.245 0.730 3.475 1.610 ;
        RECT  3.245 1.380 4.200 1.610 ;
        RECT  3.970 1.380 4.200 1.970 ;
        RECT  3.970 1.630 4.310 1.970 ;
        RECT  1.885 0.730 2.115 2.410 ;
        RECT  1.885 2.180 2.580 2.410 ;
        RECT  2.350 2.180 2.580 3.505 ;
        RECT  2.240 3.165 2.580 3.505 ;
    END
END BTHX2

MACRO BTHX16
    CLASS CORE ;
    FOREIGN BTHX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.530 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.916  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.025 2.070 6.315 2.395 ;
        RECT  5.165 2.070 5.545 2.630 ;
        RECT  5.025 2.070 5.545 2.410 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 9.697  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.970 0.700 19.405 4.150 ;
        RECT  10.325 1.840 19.405 2.440 ;
        RECT  17.530 0.700 17.870 4.150 ;
        RECT  17.520 0.700 17.870 2.440 ;
        RECT  16.090 0.700 16.435 4.150 ;
        RECT  16.080 0.700 16.435 2.440 ;
        RECT  14.650 0.700 14.990 4.150 ;
        RECT  14.645 0.700 14.990 2.440 ;
        RECT  13.210 0.700 13.550 4.150 ;
        RECT  13.205 0.700 13.550 2.440 ;
        RECT  11.855 1.840 12.195 3.415 ;
        RECT  11.770 0.700 12.120 2.440 ;
        RECT  10.585 1.840 10.925 3.415 ;
        RECT  10.325 0.700 10.665 2.440 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.255  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 3.470 1.790 4.250 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 19.530 0.400 ;
        RECT  18.250 -0.400 18.590 1.570 ;
        RECT  16.810 -0.400 17.150 1.570 ;
        RECT  15.370 -0.400 15.710 1.575 ;
        RECT  13.930 -0.400 14.270 1.570 ;
        RECT  12.490 -0.400 12.830 1.570 ;
        RECT  11.045 -0.400 11.385 1.570 ;
        RECT  9.565 -0.400 9.905 1.280 ;
        RECT  8.145 -0.400 8.485 1.510 ;
        RECT  6.705 -0.400 7.045 1.115 ;
        RECT  5.265 -0.400 5.605 1.115 ;
        RECT  2.385 -0.400 2.725 1.555 ;
        RECT  0.905 -0.400 1.245 1.650 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 19.530 5.280 ;
        RECT  18.250 2.740 18.590 5.280 ;
        RECT  16.810 2.730 17.150 5.280 ;
        RECT  15.370 2.740 15.710 5.280 ;
        RECT  13.930 2.740 14.270 5.280 ;
        RECT  12.490 3.810 12.830 5.280 ;
        RECT  11.220 3.810 11.560 5.280 ;
        RECT  9.950 3.800 10.290 5.280 ;
        RECT  8.145 3.150 8.485 5.280 ;
        RECT  6.705 3.150 7.045 5.280 ;
        RECT  5.265 3.320 5.605 5.280 ;
        RECT  2.385 3.145 2.725 5.280 ;
        RECT  0.905 2.690 1.245 3.030 ;
        RECT  0.905 2.690 1.205 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.880 1.435 2.220 ;
        RECT  0.180 0.700 0.520 4.180 ;
        RECT  3.825 1.115 4.165 1.995 ;
        RECT  3.825 1.765 4.775 1.995 ;
        RECT  4.545 1.765 4.775 4.250 ;
        RECT  1.665 2.685 3.445 2.915 ;
        RECT  5.985 2.625 9.715 2.920 ;
        RECT  4.545 2.860 6.325 3.090 ;
        RECT  1.665 2.685 2.005 3.240 ;
        RECT  3.105 2.685 3.445 4.250 ;
        RECT  5.985 2.625 6.325 4.125 ;
        RECT  7.425 2.625 7.765 4.125 ;
        RECT  8.865 2.625 9.715 4.140 ;
        RECT  4.545 2.640 4.885 4.250 ;
        RECT  3.105 4.020 4.885 4.250 ;
        RECT  3.105 0.630 4.885 0.885 ;
        RECT  4.545 0.630 4.885 1.535 ;
        RECT  5.985 0.740 6.325 1.620 ;
        RECT  4.545 1.305 5.135 1.535 ;
        RECT  8.865 0.940 9.210 1.970 ;
        RECT  4.955 1.390 7.765 1.620 ;
        RECT  7.425 0.740 7.765 1.970 ;
        RECT  7.415 1.390 7.765 1.970 ;
        RECT  8.865 1.610 10.095 1.970 ;
        RECT  7.415 1.740 10.095 1.970 ;
        RECT  1.665 1.215 2.005 2.455 ;
        RECT  3.105 0.630 3.445 2.455 ;
        RECT  9.230 1.610 9.570 2.395 ;
        RECT  1.665 2.225 4.165 2.455 ;
        RECT  3.825 2.225 4.165 3.790 ;
        RECT  5.985 2.625 8.60 2.920 ;
        RECT  4.955 1.390 6.50 1.620 ;
        RECT  7.415 1.740 9.30 1.970 ;
        RECT  1.665 2.225 3.40 2.455 ;
    END
END BTHX16

MACRO BTHX12
    CLASS CORE ;
    FOREIGN BTHX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.380 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 2.272  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.005 2.070 6.295 2.410 ;
        RECT  5.165 2.070 5.545 2.630 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.258  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  15.140 0.700 15.625 4.150 ;
        RECT  9.375 1.840 15.625 2.390 ;
        RECT  15.130 0.700 15.625 2.390 ;
        RECT  13.700 0.700 14.040 4.150 ;
        RECT  13.695 0.700 14.040 2.390 ;
        RECT  12.260 0.700 12.600 4.150 ;
        RECT  12.255 0.700 12.600 2.390 ;
        RECT  10.820 0.700 11.170 2.390 ;
        RECT  10.820 0.700 11.160 4.150 ;
        RECT  9.375 0.700 9.715 4.150 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.060  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 3.470 1.790 4.250 ;
        END
    END E
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 16.380 0.400 ;
        RECT  15.855 -0.400 16.200 1.570 ;
        RECT  14.420 -0.400 14.760 1.575 ;
        RECT  12.980 -0.400 13.320 1.570 ;
        RECT  11.540 -0.400 11.880 1.570 ;
        RECT  10.095 -0.400 10.435 1.570 ;
        RECT  8.165 -0.400 8.505 1.510 ;
        RECT  6.685 -0.400 7.025 1.115 ;
        RECT  5.245 -0.400 5.585 1.115 ;
        RECT  2.385 -0.400 2.725 1.570 ;
        RECT  0.905 -0.400 1.245 1.620 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 16.380 5.280 ;
        RECT  15.860 2.730 16.200 5.280 ;
        RECT  14.420 2.740 14.760 5.280 ;
        RECT  12.980 2.740 13.320 5.280 ;
        RECT  11.540 2.740 11.880 5.280 ;
        RECT  10.100 2.740 10.440 5.280 ;
        RECT  8.125 2.830 8.955 5.280 ;
        RECT  6.685 3.150 7.025 5.280 ;
        RECT  5.245 3.320 5.585 5.280 ;
        RECT  2.385 3.145 2.725 5.280 ;
        RECT  0.905 2.690 1.245 3.030 ;
        RECT  0.905 2.690 1.205 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.880 1.435 2.220 ;
        RECT  0.180 0.810 0.520 3.910 ;
        RECT  3.085 0.795 4.865 1.050 ;
        RECT  4.525 0.795 4.865 1.535 ;
        RECT  5.965 0.740 6.305 1.620 ;
        RECT  4.525 1.305 5.115 1.535 ;
        RECT  4.935 1.390 7.745 1.620 ;
        RECT  7.405 0.740 7.745 1.970 ;
        RECT  7.395 1.390 7.745 1.970 ;
        RECT  8.800 1.140 9.140 1.970 ;
        RECT  7.395 1.740 9.140 1.970 ;
        RECT  1.665 1.215 2.005 2.455 ;
        RECT  3.085 0.795 3.425 2.455 ;
        RECT  1.665 2.225 4.145 2.455 ;
        RECT  3.805 2.225 4.145 3.770 ;
        RECT  3.805 1.280 4.145 1.995 ;
        RECT  3.805 1.765 4.755 1.995 ;
        RECT  7.405 2.280 9.145 2.600 ;
        RECT  4.525 1.765 4.755 4.230 ;
        RECT  1.665 2.685 3.425 2.915 ;
        RECT  5.965 2.690 7.745 2.920 ;
        RECT  4.525 2.860 6.305 3.090 ;
        RECT  1.665 2.685 2.005 3.205 ;
        RECT  3.085 2.685 3.425 4.230 ;
        RECT  5.965 2.690 6.305 4.125 ;
        RECT  7.405 2.280 7.745 4.125 ;
        RECT  4.525 2.640 4.865 4.230 ;
        RECT  3.085 4.000 4.865 4.230 ;
        RECT  4.935 1.390 6.60 1.620 ;
        RECT  1.665 2.225 3.50 2.455 ;
    END
END BTHX12

MACRO BTHX1
    CLASS CORE ;
    FOREIGN BTHX1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.290 1.640 3.660 2.325 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 1.056  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 2.645 4.925 3.965 ;
        RECT  4.610 0.910 4.925 3.965 ;
        RECT  4.520 0.910 4.925 1.260 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.299  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.115 1.135 2.755 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.800 2.645 4.140 5.280 ;
        RECT  0.780 4.005 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.760 -0.400 4.100 0.710 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.545 1.595 1.885 ;
        RECT  1.365 1.545 1.595 2.985 ;
        RECT  1.365 2.640 2.110 2.985 ;
        RECT  0.180 1.025 0.520 3.545 ;
        RECT  2.380 1.115 2.720 1.950 ;
        RECT  2.380 1.720 3.060 1.950 ;
        RECT  2.830 1.720 3.060 4.075 ;
        RECT  2.830 2.750 3.300 3.090 ;
        RECT  1.540 3.245 1.880 4.075 ;
        RECT  2.830 2.750 3.115 4.075 ;
        RECT  1.540 3.735 3.115 4.075 ;
        RECT  1.880 0.635 3.310 0.865 ;
        RECT  3.080 0.635 3.310 1.410 ;
        RECT  1.880 0.635 2.115 1.315 ;
        RECT  1.580 0.975 2.115 1.315 ;
        RECT  3.080 1.110 4.290 1.410 ;
        RECT  4.040 1.110 4.290 1.970 ;
        RECT  4.040 1.630 4.380 1.970 ;
        RECT  1.885 0.635 2.115 2.410 ;
        RECT  1.885 2.180 2.600 2.410 ;
        RECT  2.370 2.180 2.600 3.505 ;
        RECT  2.260 3.165 2.600 3.505 ;
    END
END BTHX1

MACRO BTHX0
    CLASS CORE ;
    FOREIGN BTHX0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.128  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.360 2.240 4.285 2.580 ;
        END
    END A
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.480 3.340 4.915 3.680 ;
        RECT  4.600 0.910 4.915 3.680 ;
        RECT  4.480 0.910 4.915 1.410 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.256  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.820 1.135 3.800 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.680 4.080 4.020 5.280 ;
        RECT  0.780 4.120 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.815 -0.400 4.145 0.710 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.475 1.595 1.815 ;
        RECT  1.365 1.475 1.595 3.020 ;
        RECT  1.365 2.730 2.145 3.020 ;
        RECT  0.180 1.110 0.520 3.590 ;
        RECT  2.380 1.165 3.125 1.450 ;
        RECT  2.895 1.165 3.125 3.060 ;
        RECT  3.080 2.810 4.370 3.115 ;
        RECT  1.580 3.250 1.920 3.950 ;
        RECT  3.080 2.810 3.420 3.950 ;
        RECT  1.580 3.720 3.420 3.950 ;
        RECT  1.835 0.650 3.585 0.935 ;
        RECT  1.580 0.910 2.065 1.245 ;
        RECT  3.355 0.650 3.585 1.950 ;
        RECT  1.835 0.650 2.065 1.945 ;
        RECT  1.835 1.715 2.665 1.945 ;
        RECT  3.355 1.620 4.370 1.950 ;
        RECT  2.380 1.715 2.665 3.490 ;
        RECT  2.380 3.175 2.695 3.490 ;
    END
END BTHX0

MACRO BTHCX8
    CLASS CORE ;
    FOREIGN BTHCX8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.710 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 5.101  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.310 1.765 10.585 2.265 ;
        RECT  10.190 0.700 10.585 2.265 ;
        RECT  9.470 1.765 9.810 4.180 ;
        RECT  8.750 0.700 9.090 2.265 ;
        RECT  8.030 1.765 8.370 3.430 ;
        RECT  7.310 0.700 7.650 2.960 ;
        RECT  6.690 2.620 7.650 2.960 ;
        RECT  5.870 1.270 7.650 1.500 ;
        RECT  6.690 2.620 7.030 3.430 ;
        RECT  5.350 2.830 7.030 3.170 ;
        RECT  5.870 0.700 6.210 1.500 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.785  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.655 2.105 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.934  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.880 1.640 5.545 2.100 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.710 5.280 ;
        RECT  10.190 2.640 10.530 5.280 ;
        RECT  8.750 2.620 9.090 5.280 ;
        RECT  7.360 3.620 7.700 5.280 ;
        RECT  6.020 3.660 6.360 5.280 ;
        RECT  3.580 3.910 3.920 5.280 ;
        RECT  2.060 3.960 2.400 5.280 ;
        RECT  0.940 3.960 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.710 0.400 ;
        RECT  9.470 -0.400 9.810 1.535 ;
        RECT  8.030 -0.400 8.370 1.535 ;
        RECT  6.590 -0.400 6.930 1.040 ;
        RECT  5.150 -0.400 5.490 1.275 ;
        RECT  3.430 -0.400 3.770 0.710 ;
        RECT  1.415 -0.400 1.755 1.365 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.655 0.905 1.185 1.245 ;
        RECT  0.885 1.690 3.195 2.030 ;
        RECT  0.885 0.905 1.185 2.895 ;
        RECT  0.180 2.640 1.185 2.895 ;
        RECT  0.180 2.640 0.520 3.560 ;
        RECT  2.665 0.955 4.080 1.295 ;
        RECT  1.500 2.640 4.080 2.935 ;
        RECT  3.780 0.955 4.080 3.680 ;
        RECT  1.500 2.640 1.840 3.560 ;
        RECT  2.820 2.640 3.160 3.560 ;
        RECT  3.780 3.400 5.280 3.680 ;
        RECT  4.940 3.400 5.280 4.250 ;
        RECT  5.775 1.730 6.585 2.070 ;
        RECT  4.310 0.700 4.650 2.600 ;
        RECT  5.775 1.730 6.045 2.600 ;
        RECT  4.310 2.330 6.045 2.600 ;
        RECT  4.570 2.330 4.910 3.110 ;
        RECT  0.885 1.690 2.20 2.030 ;
        RECT  1.500 2.640 3.60 2.935 ;
    END
END BTHCX8

MACRO BTHCX6
    CLASS CORE ;
    FOREIGN BTHCX6 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 4.035  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.985 1.830 8.695 2.170 ;
        RECT  8.145 1.640 8.695 2.170 ;
        RECT  8.145 0.700 8.485 2.170 ;
        RECT  7.425 1.830 7.765 4.190 ;
        RECT  6.705 0.700 7.045 2.170 ;
        RECT  5.985 1.310 6.325 4.170 ;
        RECT  4.545 2.790 6.325 3.090 ;
        RECT  5.265 1.310 6.325 1.610 ;
        RECT  5.265 0.700 5.605 1.610 ;
        RECT  4.545 2.790 4.885 4.170 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.562  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.595 0.625 2.075 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.877  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.155 1.640 4.890 2.030 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  8.145 2.640 8.485 5.280 ;
        RECT  6.705 2.640 7.045 5.280 ;
        RECT  5.265 3.320 5.605 5.280 ;
        RECT  3.710 3.830 4.050 5.280 ;
        RECT  2.220 2.740 2.565 5.280 ;
        RECT  0.740 3.460 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.425 -0.400 7.765 1.580 ;
        RECT  5.985 -0.400 6.325 1.080 ;
        RECT  4.545 -0.400 4.885 1.275 ;
        RECT  2.765 -0.400 3.105 0.755 ;
        RECT  0.780 -0.400 1.120 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.025 1.155 1.365 ;
        RECT  0.855 1.625 2.580 1.965 ;
        RECT  0.855 1.025 1.155 3.020 ;
        RECT  0.180 2.680 1.155 3.020 ;
        RECT  2.050 0.985 3.140 1.325 ;
        RECT  1.500 2.210 3.140 2.510 ;
        RECT  2.840 0.985 3.140 3.600 ;
        RECT  2.840 3.260 4.290 3.600 ;
        RECT  1.500 2.210 1.840 4.180 ;
        RECT  3.430 0.935 4.025 1.275 ;
        RECT  3.430 0.935 3.775 2.560 ;
        RECT  5.120 1.840 5.460 2.560 ;
        RECT  3.430 2.260 5.460 2.560 ;
        RECT  3.430 2.260 4.40 2.560 ;
        RECT  3.430 0.935 3.770 3.030 ;
    END
END BTHCX6

MACRO BTHCX4
    CLASS CORE ;
    FOREIGN BTHCX4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 2.655  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 1.640 6.750 2.020 ;
        RECT  6.410 0.700 6.750 2.020 ;
        RECT  5.690 1.640 6.030 4.190 ;
        RECT  4.510 3.240 6.030 3.580 ;
        RECT  5.145 1.640 6.030 2.040 ;
        RECT  5.145 1.010 5.445 2.040 ;
        RECT  4.970 1.010 5.445 1.350 ;
        RECT  4.250 3.720 4.740 4.060 ;
        RECT  4.510 3.240 4.740 4.060 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.551  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.595 0.625 2.075 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.690  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.440 1.640 4.915 2.020 ;
        RECT  4.440 0.940 4.740 2.020 ;
        RECT  3.650 0.940 4.740 1.170 ;
        RECT  3.650 0.645 3.980 1.170 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 2.640 6.750 5.280 ;
        RECT  4.970 3.840 5.310 5.280 ;
        RECT  3.530 3.720 3.870 5.280 ;
        RECT  2.220 2.740 2.565 5.280 ;
        RECT  0.740 3.460 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.370 ;
        RECT  4.210 -0.400 4.550 0.710 ;
        RECT  2.765 -0.400 3.105 0.755 ;
        RECT  0.780 -0.400 1.120 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.025 1.155 1.365 ;
        RECT  0.855 1.625 2.580 1.965 ;
        RECT  0.855 1.025 1.155 3.020 ;
        RECT  0.180 2.680 1.155 3.020 ;
        RECT  3.410 1.400 3.780 2.685 ;
        RECT  3.410 2.345 4.275 2.685 ;
        RECT  3.410 1.400 3.710 2.980 ;
        RECT  2.050 0.985 3.140 1.325 ;
        RECT  1.500 2.210 3.140 2.510 ;
        RECT  2.840 0.985 3.140 3.490 ;
        RECT  3.940 3.015 4.280 3.490 ;
        RECT  2.840 3.210 4.280 3.490 ;
        RECT  1.500 2.210 1.840 4.180 ;
    END
END BTHCX4

MACRO BTHCX20
    CLASS CORE ;
    FOREIGN BTHCX20 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.900 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 12.556  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  18.380 1.810 18.720 3.520 ;
        RECT  9.010 1.810 18.720 2.480 ;
        RECT  17.650 0.700 18.145 2.480 ;
        RECT  17.080 1.810 17.420 3.520 ;
        RECT  16.210 0.700 16.550 2.480 ;
        RECT  15.780 1.810 16.120 3.520 ;
        RECT  14.770 0.700 15.110 2.480 ;
        RECT  14.480 1.810 14.820 3.515 ;
        RECT  13.330 0.700 13.670 2.480 ;
        RECT  13.180 1.810 13.520 3.520 ;
        RECT  11.890 0.700 12.230 2.480 ;
        RECT  11.880 1.810 12.220 3.520 ;
        RECT  10.580 1.810 10.920 3.520 ;
        RECT  10.450 0.700 10.790 2.480 ;
        RECT  9.280 1.810 9.620 3.520 ;
        RECT  9.010 0.700 9.350 2.795 ;
        RECT  6.745 2.410 9.620 2.795 ;
        RECT  7.570 1.340 9.350 1.570 ;
        RECT  7.980 2.410 8.320 3.520 ;
        RECT  7.570 0.700 7.910 1.570 ;
        RECT  6.745 2.410 7.085 3.520 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.451  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.510 2.460 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.531  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.395 5.585 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 18.900 5.280 ;
        RECT  17.730 3.730 18.070 5.280 ;
        RECT  16.430 3.730 16.770 5.280 ;
        RECT  15.130 3.730 15.470 5.280 ;
        RECT  13.830 3.730 14.170 5.280 ;
        RECT  12.530 3.740 12.870 5.280 ;
        RECT  11.230 3.730 11.570 5.280 ;
        RECT  9.930 3.730 10.270 5.280 ;
        RECT  8.630 3.730 8.970 5.280 ;
        RECT  7.330 3.840 7.670 5.280 ;
        RECT  4.220 3.245 4.560 5.280 ;
        RECT  2.780 3.165 3.120 5.280 ;
        RECT  0.180 3.960 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 18.900 0.400 ;
        RECT  18.375 -0.400 18.715 1.580 ;
        RECT  16.930 -0.400 17.270 1.580 ;
        RECT  15.490 -0.400 15.830 1.580 ;
        RECT  14.050 -0.400 14.390 1.580 ;
        RECT  12.610 -0.400 12.950 1.580 ;
        RECT  11.170 -0.400 11.510 1.580 ;
        RECT  9.730 -0.400 10.070 1.580 ;
        RECT  8.290 -0.400 8.630 1.110 ;
        RECT  6.850 -0.400 7.190 1.320 ;
        RECT  5.110 -0.400 5.450 1.165 ;
        RECT  3.330 -0.400 3.670 0.710 ;
        RECT  1.500 -0.400 1.840 1.460 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 1.690 3.780 2.030 ;
        RECT  0.740 1.240 1.080 3.560 ;
        RECT  2.790 1.075 3.130 1.460 ;
        RECT  2.790 1.230 4.310 1.460 ;
        RECT  4.010 1.230 4.310 3.015 ;
        RECT  2.060 2.640 4.310 2.935 ;
        RECT  3.500 2.785 5.180 3.015 ;
        RECT  4.880 2.785 5.180 4.250 ;
        RECT  6.225 2.700 6.515 4.250 ;
        RECT  2.060 2.640 2.400 4.180 ;
        RECT  3.500 2.640 3.850 4.180 ;
        RECT  6.280 2.500 6.515 4.250 ;
        RECT  4.880 3.950 6.515 4.250 ;
        RECT  4.240 0.700 4.860 1.000 ;
        RECT  5.980 0.825 6.320 2.140 ;
        RECT  5.815 1.800 8.715 2.140 ;
        RECT  4.560 0.700 4.860 2.550 ;
        RECT  5.815 1.800 6.045 2.550 ;
        RECT  4.560 2.250 6.045 2.550 ;
        RECT  5.410 2.250 5.750 3.720 ;
        RECT  0.740 1.690 2.80 2.030 ;
        RECT  2.060 2.640 3.80 2.935 ;
        RECT  5.815 1.800 7.70 2.140 ;
    END
END BTHCX20

MACRO BTHCX16
    CLASS CORE ;
    FOREIGN BTHCX16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 10.360  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  16.490 0.700 16.885 4.180 ;
        RECT  9.290 1.830 16.885 2.430 ;
        RECT  15.050 0.700 15.390 4.180 ;
        RECT  13.610 0.700 13.950 4.180 ;
        RECT  12.170 0.700 12.510 4.180 ;
        RECT  10.730 0.700 11.070 4.180 ;
        RECT  9.290 0.700 9.630 4.180 ;
        RECT  7.850 2.350 9.630 2.600 ;
        RECT  7.850 1.320 9.630 1.550 ;
        RECT  7.850 2.350 8.190 4.180 ;
        RECT  7.850 0.700 8.190 1.550 ;
        RECT  6.460 2.780 8.190 3.120 ;
        RECT  6.460 2.780 6.750 4.180 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.188  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.640 0.610 2.460 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.414  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.470 6.070 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 17.010 5.280 ;
        RECT  15.770 2.660 16.110 5.280 ;
        RECT  14.330 2.660 14.670 5.280 ;
        RECT  12.890 2.660 13.230 5.280 ;
        RECT  11.450 2.660 11.790 5.280 ;
        RECT  10.010 2.660 10.350 5.280 ;
        RECT  8.570 2.830 8.910 5.280 ;
        RECT  7.130 3.350 7.470 5.280 ;
        RECT  4.140 3.245 4.480 5.280 ;
        RECT  2.620 4.170 2.960 5.280 ;
        RECT  0.180 3.830 1.680 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 17.010 0.400 ;
        RECT  15.770 -0.400 16.110 1.600 ;
        RECT  14.330 -0.400 14.670 1.600 ;
        RECT  12.890 -0.400 13.230 1.600 ;
        RECT  11.450 -0.400 11.790 1.600 ;
        RECT  10.010 -0.400 10.350 1.600 ;
        RECT  8.570 -0.400 8.910 1.090 ;
        RECT  7.130 -0.400 7.470 1.165 ;
        RECT  5.250 -0.400 5.590 1.165 ;
        RECT  3.330 -0.400 3.670 0.710 ;
        RECT  1.560 -0.400 1.900 1.320 ;
        RECT  0.240 -0.400 0.580 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.840 1.690 3.660 2.030 ;
        RECT  0.840 1.070 1.180 3.195 ;
        RECT  0.740 2.855 1.180 3.195 ;
        RECT  2.790 1.075 3.130 1.415 ;
        RECT  2.790 1.185 4.120 1.415 ;
        RECT  3.890 1.185 4.120 3.015 ;
        RECT  2.060 2.640 4.120 2.935 ;
        RECT  3.420 2.785 5.010 3.015 ;
        RECT  2.060 2.640 2.400 3.740 ;
        RECT  4.710 2.785 5.010 4.250 ;
        RECT  3.420 2.640 3.770 4.180 ;
        RECT  5.890 2.970 6.230 4.250 ;
        RECT  4.710 3.910 6.230 4.250 ;
        RECT  4.310 0.700 4.650 1.040 ;
        RECT  6.190 0.825 6.600 1.165 ;
        RECT  6.300 1.780 8.890 2.120 ;
        RECT  4.350 0.700 4.650 2.550 ;
        RECT  6.300 0.825 6.600 2.550 ;
        RECT  4.350 2.250 6.600 2.550 ;
        RECT  5.330 2.250 5.660 3.660 ;
        RECT  0.840 1.690 2.00 2.030 ;
        RECT  2.060 2.640 3.60 2.935 ;
        RECT  6.300 1.780 7.50 2.120 ;
        RECT  4.350 2.250 5.60 2.550 ;
    END
END BTHCX16

MACRO BTHCX12
    CLASS CORE ;
    FOREIGN BTHCX12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 7.416  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  12.080 1.640 12.475 4.180 ;
        RECT  6.675 1.830 12.475 2.380 ;
        RECT  11.360 1.640 12.475 2.380 ;
        RECT  11.360 0.700 11.700 2.380 ;
        RECT  10.690 1.830 11.030 3.430 ;
        RECT  9.920 0.700 10.260 2.380 ;
        RECT  9.350 1.830 9.690 3.430 ;
        RECT  8.480 0.700 8.820 2.380 ;
        RECT  8.010 1.830 8.350 3.430 ;
        RECT  6.675 1.270 7.380 2.380 ;
        RECT  7.040 0.700 7.380 2.380 ;
        RECT  6.675 1.270 7.015 3.430 ;
        RECT  5.290 2.910 7.015 3.210 ;
        RECT  5.600 1.270 7.380 1.535 ;
        RECT  5.600 0.700 5.940 1.535 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.955  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.635 0.600 2.150 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 1.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.020 2.220 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 12.600 5.280 ;
        RECT  11.360 3.620 11.700 5.280 ;
        RECT  10.020 3.620 10.360 5.280 ;
        RECT  8.680 3.620 9.020 5.280 ;
        RECT  7.340 3.625 7.680 5.280 ;
        RECT  6.010 3.660 6.350 5.280 ;
        RECT  3.580 3.910 3.920 5.280 ;
        RECT  2.060 4.170 2.400 5.280 ;
        RECT  0.940 4.170 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 12.600 0.400 ;
        RECT  12.080 -0.400 12.420 1.310 ;
        RECT  10.640 -0.400 10.980 1.580 ;
        RECT  9.200 -0.400 9.540 1.580 ;
        RECT  7.760 -0.400 8.100 1.580 ;
        RECT  6.320 -0.400 6.660 1.040 ;
        RECT  4.880 -0.400 5.220 1.310 ;
        RECT  3.100 -0.400 3.440 0.710 ;
        RECT  1.360 -0.400 1.700 1.460 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.580 0.905 1.130 1.245 ;
        RECT  0.830 1.690 3.120 2.030 ;
        RECT  0.830 0.905 1.130 2.895 ;
        RECT  0.180 2.640 1.130 2.895 ;
        RECT  0.180 2.640 0.520 3.910 ;
        RECT  2.590 1.075 3.655 1.415 ;
        RECT  3.355 1.075 3.655 2.935 ;
        RECT  1.500 2.640 3.655 2.935 ;
        RECT  2.820 2.640 3.160 3.680 ;
        RECT  2.820 3.440 5.270 3.680 ;
        RECT  1.500 2.640 1.840 3.760 ;
        RECT  4.930 3.440 5.270 4.250 ;
        RECT  4.010 0.700 4.345 1.510 ;
        RECT  5.315 1.765 6.125 2.105 ;
        RECT  4.010 0.700 4.305 2.680 ;
        RECT  5.315 1.765 5.655 2.680 ;
        RECT  4.010 2.450 5.655 2.680 ;
        RECT  4.570 2.450 4.910 3.210 ;
        RECT  0.830 1.690 2.60 2.030 ;
        RECT  1.500 2.640 2.30 2.935 ;
        RECT  2.820 3.440 4.20 3.680 ;
    END
END BTHCX12

MACRO AO33X4
    CLASS CORE ;
    FOREIGN AO33X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.290 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.250 1.880 3.675 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.830 1.640 6.285 2.260 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.020 5.600 2.620 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.605 1.640 3.020 2.270 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 1.640 4.935 2.385 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.153  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.480 1.120 1.915 1.460 ;
        RECT  1.385 2.750 1.775 3.240 ;
        RECT  1.385 2.095 1.710 3.240 ;
        RECT  1.480 1.120 1.710 3.240 ;
        RECT  0.180 2.095 1.710 2.325 ;
        RECT  0.180 0.790 0.520 3.090 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  3.530 3.340 3.870 5.280 ;
        RECT  2.090 3.540 2.430 5.280 ;
        RECT  0.845 3.570 1.185 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.280 -0.400 6.620 0.900 ;
        RECT  2.290 -0.400 2.630 0.710 ;
        RECT  0.910 -0.400 1.250 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.810 2.860 4.590 3.110 ;
        RECT  4.250 2.860 4.590 4.160 ;
        RECT  2.810 2.860 3.150 4.160 ;
        RECT  5.685 3.320 6.030 4.160 ;
        RECT  4.250 3.890 6.030 4.160 ;
        RECT  4.295 0.630 4.635 1.410 ;
        RECT  2.145 1.130 6.750 1.410 ;
        RECT  2.145 1.130 2.375 2.285 ;
        RECT  1.955 1.945 2.375 2.285 ;
        RECT  4.970 2.850 6.750 3.080 ;
        RECT  4.970 2.850 5.310 3.660 ;
        RECT  6.515 1.130 6.750 4.160 ;
        RECT  6.410 2.850 6.750 4.160 ;
        RECT  2.145 1.130 5.40 1.410 ;
    END
END AO33X4

MACRO AO33X2
    CLASS CORE ;
    FOREIGN AO33X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.635 3.660 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.620 1.990 3.045 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.510 5.640 2.150 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.530 2.020 4.935 2.620 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.885 1.640 2.390 2.270 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 1.510 4.300 2.105 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 2.640 1.135 3.560 ;
        RECT  0.740 1.250 1.080 1.590 ;
        RECT  0.740 1.250 0.970 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  2.900 3.340 3.240 5.280 ;
        RECT  1.460 2.640 1.800 5.280 ;
        RECT  0.180 3.960 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.420 -0.400 5.760 0.710 ;
        RECT  1.550 -0.400 1.890 0.710 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.180 2.860 3.960 3.110 ;
        RECT  2.180 2.860 2.520 3.760 ;
        RECT  3.620 2.860 3.960 4.220 ;
        RECT  5.055 3.310 5.400 4.220 ;
        RECT  3.620 3.990 5.400 4.220 ;
        RECT  1.330 0.940 6.120 1.280 ;
        RECT  1.330 0.940 1.560 2.220 ;
        RECT  1.215 1.880 1.560 2.220 ;
        RECT  4.340 2.850 6.120 3.080 ;
        RECT  4.340 2.850 4.680 3.760 ;
        RECT  5.880 0.940 6.120 3.760 ;
        RECT  5.780 2.850 6.120 3.760 ;
        RECT  1.330 0.940 5.80 1.280 ;
    END
END AO33X2

MACRO AO33X1
    CLASS CORE ;
    FOREIGN AO33X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.850 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 1.510 3.030 2.150 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.395 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.510 4.965 2.070 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.020 4.305 2.620 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.640 1.760 2.170 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  2.380 3.340 2.720 5.280 ;
        RECT  0.900 2.855 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.790 -0.400 5.130 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 3.410 3.110 ;
        RECT  1.660 2.860 2.000 3.620 ;
        RECT  3.180 2.860 3.410 4.070 ;
        RECT  3.180 3.730 4.640 4.070 ;
        RECT  0.750 0.940 5.460 1.280 ;
        RECT  0.750 0.940 0.980 2.625 ;
        RECT  0.585 2.285 0.980 2.625 ;
        RECT  5.230 0.940 5.460 3.200 ;
        RECT  3.740 2.850 5.460 3.200 ;
        RECT  0.750 0.940 4.40 1.280 ;
    END
END AO33X1

MACRO AO33X0
    CLASS CORE ;
    FOREIGN AO33X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.520 3.870 ;
        RECT  0.125 0.700 0.520 1.040 ;
        RECT  0.125 0.700 0.355 3.870 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.585 2.630 ;
        RECT  2.300 1.810 2.585 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.425 1.970 2.020 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.500 3.655 2.100 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.390 4.915 2.085 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.985 1.140 2.715 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.865 2.195 4.285 2.830 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  0.980 3.530 2.265 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.520 -0.400 4.860 0.710 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.370 2.330 1.660 3.165 ;
        RECT  1.370 2.935 2.980 3.165 ;
        RECT  2.750 2.935 2.980 3.870 ;
        RECT  2.750 3.530 4.030 3.870 ;
        RECT  2.705 0.700 3.045 1.170 ;
        RECT  0.755 0.940 3.045 1.170 ;
        RECT  0.755 0.940 0.985 1.740 ;
        RECT  0.585 1.400 0.985 1.740 ;
        RECT  2.815 0.700 3.045 2.560 ;
        RECT  2.815 2.330 3.635 2.560 ;
        RECT  3.320 2.330 3.635 3.290 ;
        RECT  3.320 3.060 4.860 3.290 ;
        RECT  4.520 3.060 4.860 3.870 ;
        RECT  0.755 0.940 2.90 1.170 ;
    END
END AO33X0

MACRO AO333X1
    CLASS CORE ;
    FOREIGN AO333X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.025 4.305 2.620 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.510 1.760 2.020 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.510 4.915 2.150 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.415 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.840 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.250 6.525 2.620 ;
        END
    END H
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.510 3.030 2.105 ;
        END
    END C
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.510 6.985 2.020 ;
        END
    END G
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.510 5.885 2.020 ;
        END
    END J
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  2.380 3.320 2.720 5.280 ;
        RECT  0.900 2.840 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  4.790 -0.400 5.605 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 3.430 3.090 ;
        RECT  1.660 2.860 2.000 3.570 ;
        RECT  3.180 2.860 3.430 4.250 ;
        RECT  3.180 3.910 4.640 4.250 ;
        RECT  3.740 2.920 6.730 3.260 ;
        RECT  0.750 0.940 7.445 1.280 ;
        RECT  0.750 0.940 0.980 1.800 ;
        RECT  0.585 1.460 0.980 1.800 ;
        RECT  7.215 0.940 7.445 4.250 ;
        RECT  5.830 3.905 7.445 4.250 ;
        RECT  3.740 2.920 5.50 3.260 ;
        RECT  0.750 0.940 6.60 1.280 ;
    END
END AO333X1

MACRO AO333X0
    CLASS CORE ;
    FOREIGN AO333X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.880 0.520 4.085 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.820 1.510 4.285 2.035 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.585 1.400 3.030 1.970 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.855 2.130 2.405 2.630 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 2.200 3.655 2.630 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.500 2.120 4.970 2.645 ;
        END
    END D
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.700 1.610 6.175 2.200 ;
        END
    END H
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.950 3.470 5.555 3.900 ;
        END
    END J
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END A
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.405 1.420 6.815 2.030 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.750 -0.400 5.090 0.710 ;
        RECT  1.235 -0.400 1.575 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  0.980 3.840 2.350 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.410 2.940 3.040 3.280 ;
        RECT  2.810 2.940 3.040 4.180 ;
        RECT  2.810 3.840 4.210 4.180 ;
        RECT  3.270 2.900 5.010 3.240 ;
        RECT  3.270 2.995 6.355 3.240 ;
        RECT  6.070 2.995 6.355 3.335 ;
        RECT  3.030 0.680 3.370 1.170 ;
        RECT  6.410 0.680 6.750 1.170 ;
        RECT  0.750 0.940 6.750 1.170 ;
        RECT  0.750 0.940 1.090 1.540 ;
        RECT  5.240 0.940 5.470 2.765 ;
        RECT  5.240 2.535 6.815 2.765 ;
        RECT  6.585 2.535 6.815 4.180 ;
        RECT  5.845 3.840 6.815 4.180 ;
        RECT  3.270 2.995 5.80 3.240 ;
        RECT  0.750 0.940 5.50 1.170 ;
    END
END AO333X0

MACRO AO332X1
    CLASS CORE ;
    FOREIGN AO332X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.130 2.250 5.775 2.620 ;
        END
    END G
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.740 1.510 6.175 2.020 ;
        END
    END H
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.850 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.635 3.030 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.900 2.415 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.510 4.915 2.150 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.025 4.305 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.640 1.760 2.270 ;
        END
    END A
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.790 -0.400 5.130 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  2.380 3.320 2.720 5.280 ;
        RECT  0.900 2.855 1.240 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 3.460 3.090 ;
        RECT  1.660 2.860 2.000 3.570 ;
        RECT  3.180 2.860 3.460 4.190 ;
        RECT  3.180 3.850 4.640 4.190 ;
        RECT  0.750 0.940 6.655 1.280 ;
        RECT  0.750 0.940 0.980 2.625 ;
        RECT  0.585 2.285 0.980 2.625 ;
        RECT  6.405 0.940 6.655 3.260 ;
        RECT  5.790 2.910 6.655 3.260 ;
        RECT  3.740 2.920 5.490 3.260 ;
        RECT  5.200 2.920 5.490 4.190 ;
        RECT  5.200 3.845 6.660 4.190 ;
        RECT  0.750 0.940 5.70 1.280 ;
    END
END AO332X1

MACRO AO332X0
    CLASS CORE ;
    FOREIGN AO332X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.520 3.965 ;
        RECT  0.125 0.880 0.490 1.220 ;
        RECT  0.125 0.880 0.465 3.965 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 1.620 4.305 2.195 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.555 3.150 2.020 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 2.120 2.395 2.630 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 2.250 3.655 2.630 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.395 2.860 4.925 3.445 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.070 1.610 5.545 2.170 ;
        END
    END G
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.930 1.470 2.270 ;
        RECT  0.755 1.930 1.135 2.820 ;
        END
    END A
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.785 1.400 6.175 2.020 ;
        END
    END H
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.550 -0.400 4.890 0.710 ;
        RECT  1.035 -0.400 1.375 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  0.980 3.720 2.350 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.410 2.835 1.750 3.170 ;
        RECT  1.410 2.940 3.010 3.170 ;
        RECT  2.780 2.940 3.010 4.205 ;
        RECT  2.780 3.865 3.705 4.205 ;
        RECT  3.240 2.920 4.165 3.260 ;
        RECT  3.935 2.920 4.165 4.095 ;
        RECT  3.935 3.755 5.855 4.095 ;
        RECT  2.830 0.680 3.170 1.170 ;
        RECT  5.780 0.680 6.120 1.170 ;
        RECT  0.720 0.940 6.120 1.170 ;
        RECT  0.720 0.940 1.040 1.560 ;
        RECT  4.610 0.940 4.840 2.630 ;
        RECT  4.610 2.400 5.855 2.630 ;
        RECT  5.515 2.400 5.855 3.015 ;
        RECT  0.720 0.940 5.70 1.170 ;
    END
END AO332X0

MACRO AO331X1
    CLASS CORE ;
    FOREIGN AO331X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.020 4.305 2.620 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.640 1.760 2.270 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.510 4.915 2.150 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.415 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.840 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.140 2.200 5.650 2.620 ;
        END
    END G
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.635 3.030 2.275 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  2.380 3.320 2.720 5.280 ;
        RECT  0.900 2.840 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.790 -0.400 5.130 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 3.460 3.090 ;
        RECT  1.660 2.860 2.000 3.570 ;
        RECT  3.180 2.860 3.460 4.250 ;
        RECT  3.180 3.910 4.635 4.250 ;
        RECT  3.740 2.920 5.400 3.260 ;
        RECT  0.750 0.940 6.120 1.280 ;
        RECT  0.750 0.940 0.980 1.800 ;
        RECT  0.585 1.460 0.980 1.800 ;
        RECT  5.880 0.940 6.120 3.260 ;
        RECT  5.780 2.910 6.120 3.260 ;
        RECT  0.750 0.940 5.30 1.280 ;
    END
END AO331X1

MACRO AO331X0
    CLASS CORE ;
    FOREIGN AO331X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.408  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.470 0.520 3.870 ;
        RECT  0.115 0.880 0.520 1.220 ;
        RECT  0.115 0.880 0.345 3.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.835 1.640 4.285 2.255 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.250 3.025 2.580 ;
        RECT  2.625 1.220 2.855 2.580 ;
        RECT  2.430 1.220 2.855 1.520 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.750 2.395 2.580 ;
        RECT  1.755 1.750 2.395 2.090 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.085 1.555 3.605 2.025 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.155 3.250 5.555 3.860 ;
        END
    END G
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.730 2.175 1.135 2.785 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 1.580 5.030 2.075 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.350 -0.400 4.690 0.710 ;
        RECT  1.035 -0.400 1.375 1.020 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  0.980 3.530 2.250 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.365 2.495 1.650 3.040 ;
        RECT  1.365 2.810 2.900 3.040 ;
        RECT  2.670 2.810 2.900 3.870 ;
        RECT  2.670 3.530 3.685 3.870 ;
        RECT  3.140 2.785 4.880 3.070 ;
        RECT  4.540 2.785 4.880 3.875 ;
        RECT  1.970 0.680 3.315 0.965 ;
        RECT  5.150 0.670 5.490 1.180 ;
        RECT  3.085 0.940 5.490 1.180 ;
        RECT  0.750 1.290 2.200 1.520 ;
        RECT  1.970 0.680 2.200 1.520 ;
        RECT  0.575 1.520 0.980 1.860 ;
        RECT  5.260 0.670 5.490 3.020 ;
        RECT  5.150 2.705 5.490 3.020 ;
        RECT  3.085 0.940 4.20 1.180 ;
    END
END AO331X0

MACRO AO32X4
    CLASS CORE ;
    FOREIGN AO32X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.635 4.290 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.250 1.880 3.675 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.160 2.075 5.680 2.620 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.515 1.640 3.020 2.270 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 1.510 4.930 2.195 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.180 1.360 1.825 1.700 ;
        RECT  0.180 2.920 1.800 3.260 ;
        RECT  0.755 1.360 1.135 3.260 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  3.620 3.340 3.960 5.280 ;
        RECT  2.180 2.640 2.520 5.280 ;
        RECT  0.840 3.560 1.180 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.620 -0.400 5.960 0.710 ;
        RECT  2.235 -0.400 2.575 0.710 ;
        RECT  0.865 -0.400 1.205 1.130 ;
        RECT  0.115 -0.400 1.205 0.405 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.900 2.860 4.680 3.110 ;
        RECT  4.340 2.860 4.680 4.250 ;
        RECT  2.900 2.860 3.240 4.160 ;
        RECT  5.780 3.310 6.120 4.250 ;
        RECT  4.340 4.020 6.120 4.250 ;
        RECT  2.055 0.940 6.140 1.280 ;
        RECT  2.055 0.940 2.285 2.285 ;
        RECT  1.685 1.945 2.285 2.285 ;
        RECT  5.910 0.940 6.140 3.080 ;
        RECT  5.060 2.850 6.140 3.080 ;
        RECT  5.060 2.850 5.400 3.790 ;
        RECT  2.055 0.940 5.60 1.280 ;
    END
END AO32X4

MACRO AO32X2
    CLASS CORE ;
    FOREIGN AO32X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.635 3.660 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.620 1.880 3.045 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.530 2.075 5.050 2.630 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.885 1.640 2.390 2.270 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 1.510 4.300 2.105 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.900  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.750 1.135 3.560 ;
        RECT  0.755 1.250 1.135 1.590 ;
        RECT  0.755 1.250 0.985 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  2.990 3.320 3.330 5.280 ;
        RECT  1.550 2.640 1.890 5.280 ;
        RECT  0.230 3.960 0.570 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.990 -0.400 5.330 0.710 ;
        RECT  1.605 -0.400 1.945 0.710 ;
        RECT  0.230 -0.400 0.570 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.270 2.860 4.050 3.090 ;
        RECT  2.270 2.860 2.610 3.760 ;
        RECT  3.710 2.860 4.050 4.250 ;
        RECT  5.150 3.320 5.490 4.250 ;
        RECT  3.710 4.020 5.490 4.250 ;
        RECT  1.380 0.940 5.510 1.280 ;
        RECT  1.380 0.940 1.610 2.285 ;
        RECT  1.215 1.945 1.610 2.285 ;
        RECT  5.280 0.940 5.510 3.090 ;
        RECT  4.430 2.860 5.510 3.090 ;
        RECT  4.430 2.860 4.770 3.760 ;
        RECT  1.380 0.940 4.80 1.280 ;
    END
END AO32X2

MACRO AO32X1
    CLASS CORE ;
    FOREIGN AO32X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.850 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.635 3.030 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.415 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.075 4.325 2.620 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.640 1.760 2.270 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  2.380 3.340 2.720 5.280 ;
        RECT  0.900 2.855 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.360 -0.400 4.700 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 3.410 3.110 ;
        RECT  1.660 2.860 2.000 3.635 ;
        RECT  3.180 2.860 3.410 4.070 ;
        RECT  3.180 3.730 4.640 4.070 ;
        RECT  0.750 0.940 4.785 1.280 ;
        RECT  0.750 0.940 0.980 2.625 ;
        RECT  0.585 2.285 0.980 2.625 ;
        RECT  4.555 0.940 4.785 3.200 ;
        RECT  3.740 2.850 4.785 3.200 ;
        RECT  0.750 0.940 3.90 1.280 ;
    END
END AO32X1

MACRO AO32X0
    CLASS CORE ;
    FOREIGN AO32X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.493  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.880 0.520 3.975 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.250 3.025 2.020 ;
        RECT  2.360 1.250 3.025 1.585 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.855 2.130 2.405 2.630 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 2.050 3.655 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.785 3.430 4.285 3.955 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  0.980 3.730 2.350 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.870 -0.400 4.210 1.020 ;
        RECT  0.980 -0.400 1.320 0.990 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.410 2.860 1.750 3.200 ;
        RECT  1.410 2.970 3.070 3.200 ;
        RECT  2.840 2.970 3.070 4.070 ;
        RECT  2.840 3.730 3.180 4.070 ;
        RECT  1.550 0.680 3.490 1.020 ;
        RECT  3.260 0.680 3.490 1.510 ;
        RECT  3.260 1.270 4.115 1.510 ;
        RECT  1.550 0.680 1.780 1.560 ;
        RECT  0.750 1.220 1.780 1.560 ;
        RECT  3.885 1.270 4.115 3.200 ;
        RECT  3.410 2.860 4.115 3.200 ;
    END
END AO32X0

MACRO AO322X1
    CLASS CORE ;
    FOREIGN AO322X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 2.075 4.350 2.620 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.295 1.640 1.760 2.270 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.415 2.630 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.830 0.560 1.170 ;
        RECT  0.125 2.850 0.520 3.740 ;
        RECT  0.125 0.830 0.355 3.740 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.630 1.510 6.175 2.020 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 2.250 6.000 2.620 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.635 3.030 2.275 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  2.365 3.340 2.740 5.280 ;
        RECT  0.900 2.855 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.360 -0.400 5.170 0.710 ;
        RECT  1.015 -0.400 1.355 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 3.480 3.110 ;
        RECT  1.660 2.860 2.000 3.585 ;
        RECT  3.140 2.860 3.480 4.160 ;
        RECT  3.140 3.820 4.640 4.160 ;
        RECT  3.740 2.850 5.490 3.200 ;
        RECT  5.200 2.850 5.490 4.250 ;
        RECT  5.200 3.905 6.660 4.250 ;
        RECT  0.790 0.940 6.705 1.280 ;
        RECT  0.790 0.940 1.020 2.625 ;
        RECT  0.585 2.285 1.020 2.625 ;
        RECT  6.405 0.940 6.705 3.280 ;
        RECT  5.790 2.930 6.705 3.280 ;
        RECT  0.790 0.940 5.50 1.280 ;
    END
END AO322X1

MACRO AO322X0
    CLASS CORE ;
    FOREIGN AO322X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.880 0.520 3.965 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 3.470 4.250 4.100 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.520 3.030 2.020 ;
        RECT  2.530 1.520 3.030 1.925 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.800 2.120 2.395 2.630 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.630 3.680 2.215 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.440 1.630 4.920 2.170 ;
        END
    END F
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.930 1.470 2.270 ;
        RECT  0.755 1.930 1.135 2.630 ;
        END
    END A
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.099  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.155 1.400 5.545 2.070 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.920 -0.400 4.260 0.710 ;
        RECT  1.030 -0.400 1.370 0.710 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  0.980 3.720 2.350 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  1.410 2.860 1.750 3.200 ;
        RECT  1.410 2.970 3.040 3.200 ;
        RECT  2.810 2.970 3.040 4.060 ;
        RECT  2.810 3.720 3.660 4.060 ;
        RECT  3.410 2.895 3.750 3.235 ;
        RECT  3.410 3.005 4.710 3.235 ;
        RECT  4.480 3.005 4.710 4.060 ;
        RECT  4.480 3.720 4.990 4.060 ;
        RECT  2.690 0.680 3.030 1.170 ;
        RECT  5.150 0.680 5.490 1.170 ;
        RECT  0.750 0.940 5.490 1.170 ;
        RECT  0.750 0.940 1.040 1.560 ;
        RECT  3.980 0.940 4.210 2.775 ;
        RECT  3.980 2.545 5.225 2.775 ;
        RECT  4.940 2.545 5.225 2.980 ;
        RECT  0.750 0.940 4.60 1.170 ;
    END
END AO322X0

MACRO AO321X4
    CLASS CORE ;
    FOREIGN AO321X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.489  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.270 2.335 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.715 2.250 4.235 2.630 ;
        RECT  3.715 2.195 4.075 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.045 1.640 3.655 1.970 ;
        RECT  3.045 1.640 3.385 2.460 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 1.950 5.565 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.440 1.640 4.915 2.140 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.485  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.425 2.120 2.715 2.635 ;
        RECT  2.015 2.860 2.435 3.240 ;
        RECT  2.205 2.405 2.435 3.240 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.991  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.180 1.360 1.735 1.700 ;
        RECT  0.180 2.920 1.680 3.260 ;
        RECT  0.755 1.360 1.135 3.260 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.495 -0.400 5.835 0.940 ;
        RECT  2.230 -0.400 2.570 0.950 ;
        RECT  0.815 -0.400 1.155 1.130 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  3.380 3.580 3.720 5.280 ;
        RECT  2.080 3.555 2.420 5.280 ;
        RECT  0.760 3.560 1.100 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.805 2.860 5.480 3.200 ;
        RECT  4.565 3.580 6.175 3.920 ;
        RECT  4.040 0.630 4.380 1.410 ;
        RECT  4.040 1.170 6.805 1.410 ;
        RECT  6.410 0.700 6.805 1.410 ;
        RECT  1.965 1.180 6.805 1.410 ;
        RECT  1.965 1.180 2.195 2.160 ;
        RECT  1.690 1.930 2.015 2.270 ;
        RECT  6.575 0.700 6.805 3.200 ;
        RECT  6.410 2.860 6.805 3.200 ;
        RECT  2.805 2.860 4.70 3.200 ;
        RECT  4.040 1.170 5.60 1.410 ;
        RECT  1.965 1.180 5.90 1.410 ;
    END
END AO321X4

MACRO AO321X2
    CLASS CORE ;
    FOREIGN AO321X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.640 2.310 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.350 1.120 1.175 1.430 ;
        RECT  0.755 2.640 1.155 3.560 ;
        RECT  0.350 2.640 1.155 2.870 ;
        RECT  0.350 1.120 0.585 2.870 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.985 2.250 3.685 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.415 1.640 3.025 2.020 ;
        RECT  2.415 1.640 2.755 2.460 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 2.025 4.935 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.645 1.640 4.285 2.020 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.376  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.120 2.085 2.460 ;
        RECT  1.385 2.120 1.765 3.240 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.845 -0.400 5.185 0.950 ;
        RECT  1.600 -0.400 1.940 0.950 ;
        RECT  0.275 -0.400 0.615 0.720 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  2.750 3.580 3.090 5.280 ;
        RECT  1.600 3.580 1.940 5.280 ;
        RECT  0.275 3.960 0.615 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.175 2.860 4.850 3.200 ;
        RECT  3.935 3.580 5.545 3.920 ;
        RECT  3.350 0.865 3.690 1.410 ;
        RECT  5.780 0.865 6.175 1.410 ;
        RECT  1.410 1.180 6.175 1.410 ;
        RECT  1.410 1.180 1.640 1.890 ;
        RECT  0.815 1.660 1.640 1.890 ;
        RECT  0.815 1.660 1.155 2.285 ;
        RECT  5.945 0.865 6.175 3.200 ;
        RECT  5.780 2.860 6.175 3.200 ;
        RECT  2.175 2.860 3.70 3.200 ;
        RECT  1.410 1.180 5.60 1.410 ;
    END
END AO321X2

MACRO AO321X1
    CLASS CORE ;
    FOREIGN AO321X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.510 5.080 2.020 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.840 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.510 3.030 2.105 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.415 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.510 4.305 2.105 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 1.510 3.670 2.105 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.640 1.760 2.270 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  2.380 3.340 2.720 5.280 ;
        RECT  0.900 2.840 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.350 -0.400 4.690 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.860 4.805 3.110 ;
        RECT  4.465 2.455 4.805 3.205 ;
        RECT  3.140 2.860 4.805 3.205 ;
        RECT  1.660 2.860 2.000 3.570 ;
        RECT  0.750 0.940 5.555 1.280 ;
        RECT  0.750 0.940 0.980 1.800 ;
        RECT  0.585 1.460 0.980 1.800 ;
        RECT  5.325 0.940 5.555 3.990 ;
        RECT  4.895 3.645 5.555 3.990 ;
        RECT  1.660 2.860 3.70 3.110 ;
        RECT  0.750 0.940 4.60 1.280 ;
    END
END AO321X1

MACRO AO321X0
    CLASS CORE ;
    FOREIGN AO321X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.426  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.520 4.135 ;
        RECT  0.125 0.880 0.520 1.220 ;
        RECT  0.125 0.880 0.355 4.135 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 1.640 3.025 2.420 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.585 2.405 2.185 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.025 3.675 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.305 2.450 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.480 4.925 2.030 ;
        END
    END F
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.275 1.640 1.765 2.265 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  0.980 3.890 2.395 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.720 -0.400 4.060 0.710 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.410 2.860 4.595 3.200 ;
        RECT  2.690 0.680 3.030 1.250 ;
        RECT  4.520 0.910 4.860 1.250 ;
        RECT  0.755 1.020 4.860 1.250 ;
        RECT  0.605 1.675 0.985 2.015 ;
        RECT  0.755 1.020 0.985 3.660 ;
        RECT  0.755 3.430 4.750 3.660 ;
        RECT  4.520 3.430 4.750 4.230 ;
        RECT  4.520 3.890 4.860 4.230 ;
        RECT  1.410 2.860 3.80 3.200 ;
        RECT  0.755 1.020 3.30 1.250 ;
        RECT  0.755 3.430 3.40 3.660 ;
    END
END AO321X0

MACRO AO31X4
    CLASS CORE ;
    FOREIGN AO31X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.209  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.165 1.485 1.955 1.715 ;
        RECT  1.625 0.890 1.955 1.715 ;
        RECT  0.165 2.810 1.860 3.260 ;
        RECT  0.165 0.890 0.525 1.715 ;
        RECT  0.165 0.890 0.505 3.260 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.040 1.625 5.545 2.170 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.250 2.065 3.675 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.630 3.020 2.280 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.635 4.350 2.170 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.640 3.320 3.980 5.280 ;
        RECT  2.200 3.555 2.540 5.280 ;
        RECT  0.845 3.560 1.185 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.090 -0.400 5.430 0.710 ;
        RECT  2.385 -0.400 5.430 0.405 ;
        RECT  2.385 -0.400 2.725 0.710 ;
        RECT  0.905 -0.400 1.245 1.230 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.920 2.860 4.740 3.090 ;
        RECT  2.920 2.860 3.260 4.180 ;
        RECT  4.400 2.860 4.740 4.185 ;
        RECT  2.185 0.940 4.810 1.280 ;
        RECT  2.185 0.940 2.415 2.295 ;
        RECT  1.645 1.945 2.415 2.295 ;
        RECT  4.580 0.940 4.810 2.630 ;
        RECT  4.580 2.400 5.460 2.630 ;
        RECT  5.120 2.400 5.460 4.185 ;
        RECT  2.185 0.940 3.60 1.280 ;
    END
END AO31X4

MACRO AO31X2
    CLASS CORE ;
    FOREIGN AO31X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.901  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.860 1.190 3.760 ;
        RECT  0.755 1.250 1.185 1.590 ;
        RECT  0.755 1.250 0.985 3.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.350 1.560 4.915 2.055 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.980 3.045 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.885 1.640 2.395 2.270 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.635 3.660 2.365 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.010 3.340 3.350 5.280 ;
        RECT  1.570 2.855 1.910 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.090 -0.400 4.430 0.710 ;
        RECT  1.605 -0.400 1.945 0.710 ;
        RECT  0.180 -0.400 0.520 0.720 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.290 2.860 4.110 3.110 ;
        RECT  2.290 2.860 2.630 3.760 ;
        RECT  3.770 2.860 4.110 3.760 ;
        RECT  1.415 0.940 4.120 1.280 ;
        RECT  3.890 0.940 4.120 2.630 ;
        RECT  1.415 0.940 1.645 2.480 ;
        RECT  1.215 2.140 1.645 2.480 ;
        RECT  3.890 2.400 4.830 2.630 ;
        RECT  4.490 2.400 4.830 3.760 ;
        RECT  1.415 0.940 3.70 1.280 ;
    END
END AO31X2

MACRO AO31X1
    CLASS CORE ;
    FOREIGN AO31X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.850 0.520 3.760 ;
        RECT  0.125 0.830 0.520 1.170 ;
        RECT  0.125 0.830 0.355 3.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.720 1.470 4.285 2.030 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.990 1.880 2.415 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.255 1.640 1.760 2.270 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.203  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.635 3.030 2.275 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  2.380 3.370 2.720 5.280 ;
        RECT  0.900 2.855 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.460 -0.400 3.800 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.660 2.890 3.480 3.140 ;
        RECT  3.140 2.890 3.480 3.230 ;
        RECT  1.660 2.890 2.000 3.620 ;
        RECT  0.750 0.940 3.490 1.280 ;
        RECT  3.260 0.940 3.490 2.630 ;
        RECT  0.750 0.940 0.980 2.625 ;
        RECT  0.585 2.285 0.980 2.625 ;
        RECT  3.260 2.400 4.200 2.630 ;
        RECT  3.860 2.400 4.200 3.315 ;
        RECT  0.750 0.940 2.60 1.280 ;
    END
END AO31X1

MACRO AO31X0
    CLASS CORE ;
    FOREIGN AO31X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.520 4.175 ;
        RECT  0.125 0.880 0.520 1.220 ;
        RECT  0.125 0.880 0.465 4.175 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.635 3.030 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.880 2.415 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.440 3.655 2.150 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.260 1.640 1.765 2.270 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  0.980 3.930 2.350 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.260 -0.400 3.600 0.710 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.755 0.990 2.980 1.330 ;
        RECT  0.695 1.400 0.985 1.740 ;
        RECT  0.755 0.990 0.985 3.700 ;
        RECT  0.755 3.470 3.245 3.700 ;
        RECT  2.905 3.470 3.245 4.250 ;
        RECT  1.410 2.860 3.250 3.200 ;
        RECT  0.755 0.990 1.60 1.330 ;
        RECT  0.755 3.470 2.90 3.700 ;
    END
END AO31X0

MACRO AO311X4
    CLASS CORE ;
    FOREIGN AO311X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 1.640 3.025 2.270 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.300 5.725 2.630 ;
        RECT  5.440 1.800 5.725 2.630 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.635 4.300 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 2.000 3.675 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.468  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.530 1.510 5.080 2.085 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.585 2.660 1.960 3.915 ;
        RECT  1.585 0.890 1.905 1.700 ;
        RECT  1.585 0.890 1.815 3.915 ;
        RECT  0.180 2.250 1.815 2.630 ;
        RECT  0.180 0.890 0.520 3.915 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  3.820 3.350 4.160 5.280 ;
        RECT  2.370 2.770 2.710 5.280 ;
        RECT  0.900 2.860 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.020 -0.400 5.360 0.710 ;
        RECT  2.380 -0.400 2.720 0.710 ;
        RECT  0.900 -0.400 1.240 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.090 2.860 4.880 3.120 ;
        RECT  4.540 2.860 4.880 4.180 ;
        RECT  3.090 2.860 3.430 4.185 ;
        RECT  2.135 0.940 6.185 1.280 ;
        RECT  2.135 0.940 2.365 2.305 ;
        RECT  2.045 1.950 2.365 2.305 ;
        RECT  5.955 0.940 6.185 3.090 ;
        RECT  5.695 2.860 6.035 4.180 ;
        RECT  2.135 0.940 5.70 1.280 ;
    END
END AO311X4

MACRO AO311X2
    CLASS CORE ;
    FOREIGN AO311X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.935 1.640 2.390 2.270 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.485 2.250 5.090 2.630 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.635 3.670 2.275 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.620 1.880 3.045 2.630 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 1.510 4.420 2.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 2.840 1.240 3.760 ;
        RECT  0.860 0.910 1.185 1.250 ;
        RECT  0.860 0.910 1.090 3.240 ;
        RECT  0.755 2.840 1.240 3.240 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.105 3.340 3.445 5.280 ;
        RECT  1.655 2.840 2.000 5.280 ;
        RECT  0.180 2.840 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.360 -0.400 4.700 0.710 ;
        RECT  1.660 -0.400 2.000 0.710 ;
        RECT  0.180 -0.400 0.520 1.240 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.385 2.860 4.205 3.110 ;
        RECT  2.385 2.860 2.725 3.960 ;
        RECT  3.855 2.860 4.205 3.960 ;
        RECT  1.415 0.940 5.550 1.280 ;
        RECT  1.415 0.940 1.645 2.290 ;
        RECT  1.320 1.950 1.645 2.290 ;
        RECT  5.320 0.940 5.550 3.090 ;
        RECT  5.020 2.860 5.360 3.960 ;
        RECT  1.415 0.940 4.00 1.280 ;
    END
END AO311X2

MACRO AO311X1
    CLASS CORE ;
    FOREIGN AO311X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.180 1.640 1.775 2.050 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.000 4.285 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.820  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.520 3.860 ;
        RECT  0.125 3.050 0.490 3.860 ;
        RECT  0.125 1.080 0.490 1.420 ;
        RECT  0.125 1.080 0.355 3.860 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.575 2.245 3.030 2.785 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.735 2.445 2.345 2.785 ;
        RECT  2.015 2.250 2.345 2.785 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 1.640 3.655 2.100 ;
        RECT  3.050 1.640 3.655 2.015 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  0.940 4.170 2.440 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.065 -0.400 3.405 0.710 ;
        RECT  0.975 -0.400 1.315 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.500 3.475 3.240 3.760 ;
        RECT  2.900 3.475 3.240 4.250 ;
        RECT  3.865 0.750 4.205 1.380 ;
        RECT  0.720 1.150 4.205 1.380 ;
        RECT  2.505 1.150 2.845 1.490 ;
        RECT  0.585 2.375 0.950 2.715 ;
        RECT  0.720 1.150 0.950 3.245 ;
        RECT  3.890 2.905 4.230 3.245 ;
        RECT  0.720 3.015 4.230 3.245 ;
        RECT  0.720 1.150 3.30 1.380 ;
        RECT  0.720 3.015 3.20 3.245 ;
    END
END AO311X1

MACRO AO311X0
    CLASS CORE ;
    FOREIGN AO311X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.730 0.520 4.070 ;
        RECT  0.125 0.880 0.520 1.360 ;
        RECT  0.125 0.880 0.480 1.390 ;
        RECT  0.125 0.880 0.355 4.070 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.025 2.465 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.955 2.130 2.415 2.580 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.970 3.670 2.580 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.215 1.640 1.725 2.020 ;
        RECT  1.215 1.640 1.525 2.470 ;
        END
    END A
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.900 1.540 4.285 2.175 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  0.980 3.730 2.350 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.190 -0.400 3.530 0.710 ;
        RECT  0.980 -0.400 1.320 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.410 2.755 1.750 3.040 ;
        RECT  1.410 2.810 3.250 3.040 ;
        RECT  2.490 0.970 2.830 1.310 ;
        RECT  3.890 0.970 4.230 1.310 ;
        RECT  0.755 1.080 4.230 1.310 ;
        RECT  0.585 1.595 0.985 1.935 ;
        RECT  0.755 1.080 0.985 3.500 ;
        RECT  0.755 3.270 4.050 3.500 ;
        RECT  3.710 3.270 4.050 4.070 ;
        RECT  0.755 1.080 3.70 1.310 ;
        RECT  0.755 3.270 3.70 3.500 ;
    END
END AO311X0

MACRO AO22X4
    CLASS CORE ;
    FOREIGN AO22X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 1.525 1.765 2.105 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.595 1.930 1.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.960 2.395 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.234  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.765 0.950 6.105 3.450 ;
        RECT  4.435 1.640 6.105 2.020 ;
        RECT  4.325 2.640 4.665 3.450 ;
        RECT  4.435 0.950 4.665 3.450 ;
        RECT  4.325 0.950 4.665 1.290 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.085 2.100 3.655 2.720 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.045 2.640 5.385 5.280 ;
        RECT  3.600 4.170 3.940 5.280 ;
        RECT  0.900 3.410 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.045 -0.400 5.385 1.290 ;
        RECT  2.915 -0.400 3.905 1.270 ;
        RECT  0.320 -0.400 0.660 1.280 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.885 1.960 3.180 ;
        RECT  1.620 2.885 1.960 3.825 ;
        RECT  3.085 2.950 3.400 3.825 ;
        RECT  1.620 3.595 3.400 3.825 ;
        RECT  0.180 2.885 0.520 4.180 ;
        RECT  1.600 0.945 2.275 1.285 ;
        RECT  2.045 0.945 2.275 1.730 ;
        RECT  2.045 1.500 4.205 1.730 ;
        RECT  3.885 1.500 4.205 2.040 ;
        RECT  2.625 1.500 2.855 3.365 ;
        RECT  2.340 3.025 2.855 3.365 ;
        RECT  2.045 1.500 3.60 1.730 ;
    END
END AO22X4

MACRO AO22X2
    CLASS CORE ;
    FOREIGN AO22X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.365 1.525 1.765 2.105 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.595 1.930 1.135 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.920 2.395 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.325 1.640 4.915 2.020 ;
        RECT  4.325 0.830 4.665 3.560 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.085 2.170 3.655 2.720 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.045 2.640 5.385 5.280 ;
        RECT  3.765 3.960 4.105 5.280 ;
        RECT  0.900 3.345 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.085 -0.400 5.425 1.280 ;
        RECT  2.915 -0.400 3.905 1.230 ;
        RECT  0.320 -0.400 0.660 1.200 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.885 1.960 3.115 ;
        RECT  1.620 2.885 1.960 3.995 ;
        RECT  0.180 2.885 0.520 3.995 ;
        RECT  3.085 2.950 3.400 3.995 ;
        RECT  1.620 3.765 3.400 3.995 ;
        RECT  1.600 0.850 2.275 1.190 ;
        RECT  2.045 0.850 2.275 1.690 ;
        RECT  2.045 1.460 4.095 1.690 ;
        RECT  3.755 1.460 4.095 1.800 ;
        RECT  2.625 1.460 2.855 3.535 ;
        RECT  2.340 3.195 2.855 3.535 ;
        RECT  2.045 1.460 3.50 1.690 ;
    END
END AO22X2

MACRO AO22X1
    CLASS CORE ;
    FOREIGN AO22X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.734  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 2.250 4.285 2.980 ;
        RECT  3.980 0.870 4.285 2.980 ;
        RECT  3.890 0.870 4.285 1.210 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.201  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.635 1.190 2.270 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.201  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.135 0.525 2.730 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.201  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.880 2.120 2.395 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.201  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.615 3.070 2.165 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.330 3.280 3.670 5.280 ;
        RECT  0.910 4.170 1.250 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.080 -0.400 3.420 0.885 ;
        RECT  0.180 -0.400 0.520 1.280 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 3.695 2.970 3.930 ;
        RECT  1.510 3.695 2.970 4.035 ;
        RECT  0.180 3.695 0.520 4.250 ;
        RECT  1.420 0.960 1.825 1.345 ;
        RECT  1.420 1.115 3.660 1.345 ;
        RECT  3.410 1.115 3.660 1.985 ;
        RECT  3.410 1.645 3.750 1.985 ;
        RECT  1.420 0.960 1.650 3.225 ;
        RECT  1.420 2.885 2.410 3.225 ;
        RECT  0.180 3.695 1.80 3.930 ;
        RECT  1.420 1.115 2.20 1.345 ;
    END
END AO22X1

MACRO AO22X0
    CLASS CORE ;
    FOREIGN AO22X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.453  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.470 0.520 4.175 ;
        RECT  0.125 0.880 0.520 1.220 ;
        RECT  0.125 0.880 0.355 4.175 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.122  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 1.640 2.395 2.220 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.122  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.225 2.125 1.765 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.122  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.045 3.025 2.670 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.122  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.155 3.470 3.655 4.080 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  0.980 3.655 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.260 -0.400 3.600 0.710 ;
        RECT  0.980 -0.400 1.320 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 2.860 2.410 3.200 ;
        RECT  2.180 2.860 2.410 4.250 ;
        RECT  2.180 3.930 2.520 4.250 ;
        RECT  2.230 0.910 2.570 1.410 ;
        RECT  0.750 1.180 3.485 1.410 ;
        RECT  0.750 1.180 1.090 1.560 ;
        RECT  3.255 1.180 3.485 3.240 ;
        RECT  2.780 2.900 3.485 3.240 ;
        RECT  0.750 1.180 2.30 1.410 ;
    END
END AO22X0

MACRO AO222X4
    CLASS CORE ;
    FOREIGN AO222X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 2.120 3.045 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.605 1.915 2.150 2.255 ;
        RECT  1.605 1.030 1.865 2.255 ;
        RECT  1.385 1.030 1.865 1.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.375 2.260 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.020 0.515 1.630 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.250 4.485 2.635 ;
        RECT  4.065 2.120 4.485 2.635 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.730 3.825 2.030 ;
        RECT  3.275 1.730 3.665 2.635 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.000  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.880 2.920 7.380 3.260 ;
        RECT  5.770 1.360 7.380 1.695 ;
        RECT  6.425 1.360 6.805 3.260 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.460 3.560 6.800 5.280 ;
        RECT  5.225 3.555 5.565 5.280 ;
        RECT  1.620 3.840 1.960 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.405 -0.400 6.745 1.130 ;
        RECT  5.135 -0.400 5.475 1.135 ;
        RECT  3.285 -0.400 3.625 1.040 ;
        RECT  0.810 -0.400 1.150 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 3.325 2.700 3.555 ;
        RECT  0.900 3.325 1.240 4.180 ;
        RECT  2.360 3.325 2.700 4.180 ;
        RECT  0.180 2.865 3.420 3.095 ;
        RECT  3.080 2.865 3.420 4.160 ;
        RECT  0.180 2.865 0.520 4.160 ;
        RECT  4.520 3.345 4.860 4.160 ;
        RECT  3.080 3.905 4.860 4.160 ;
        RECT  2.095 0.730 2.435 1.500 ;
        RECT  4.435 0.845 4.775 1.500 ;
        RECT  2.095 1.270 4.945 1.500 ;
        RECT  4.715 1.945 5.870 2.285 ;
        RECT  4.715 1.270 4.945 3.095 ;
        RECT  3.800 2.865 4.945 3.095 ;
        RECT  3.800 2.865 4.140 3.675 ;
        RECT  0.180 2.865 2.20 3.095 ;
        RECT  2.095 1.270 3.50 1.500 ;
    END
END AO222X4

MACRO AO222X2
    CLASS CORE ;
    FOREIGN AO222X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 2.750 6.175 3.560 ;
        RECT  5.890 1.250 6.175 3.560 ;
        RECT  5.780 1.250 6.175 1.590 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.490 2.120 3.065 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.605 1.915 2.220 2.255 ;
        RECT  1.605 1.030 1.870 2.255 ;
        RECT  1.385 1.030 1.870 1.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.375 2.230 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.020 0.515 1.630 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.195 4.475 2.635 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.295 1.610 3.825 1.950 ;
        RECT  3.295 1.610 3.665 2.635 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.340 3.960 6.680 5.280 ;
        RECT  5.220 3.960 5.560 5.280 ;
        RECT  1.620 3.840 1.960 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.340 -0.400 6.680 0.720 ;
        RECT  5.220 -0.400 5.560 0.720 ;
        RECT  3.330 -0.400 3.670 0.905 ;
        RECT  0.810 -0.400 1.150 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 3.325 2.700 3.555 ;
        RECT  0.900 3.325 1.240 4.180 ;
        RECT  2.360 3.325 2.700 4.180 ;
        RECT  0.180 2.865 3.420 3.095 ;
        RECT  3.080 2.865 3.420 4.160 ;
        RECT  0.180 2.865 0.520 4.160 ;
        RECT  4.520 3.345 4.860 4.160 ;
        RECT  3.080 3.930 4.860 4.160 ;
        RECT  2.100 0.880 2.440 1.365 ;
        RECT  4.495 0.845 4.935 1.365 ;
        RECT  2.100 1.135 4.935 1.365 ;
        RECT  4.705 1.945 5.640 2.285 ;
        RECT  4.705 0.845 4.935 3.095 ;
        RECT  3.800 2.865 4.935 3.095 ;
        RECT  3.800 2.865 4.140 3.700 ;
        RECT  0.180 2.865 2.10 3.095 ;
        RECT  2.100 1.135 3.40 1.365 ;
    END
END AO222X2

MACRO AO222X1
    CLASS CORE ;
    FOREIGN AO222X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.850 0.575 1.190 ;
        RECT  0.125 3.260 0.520 4.180 ;
        RECT  0.125 0.850 0.410 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.765 2.630 ;
        RECT  3.420 2.045 3.765 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.890 2.415 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 1.630 1.775 2.240 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.590 3.190 2.035 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.455 1.640 4.915 2.170 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.090 2.790 5.555 3.315 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  0.900 2.860 2.040 3.150 ;
        RECT  0.900 2.860 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.760 -0.400 4.100 0.860 ;
        RECT  1.055 -0.400 1.395 0.860 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.420 2.860 4.080 3.145 ;
        RECT  2.420 2.860 2.650 4.060 ;
        RECT  1.660 3.720 2.650 4.060 ;
        RECT  3.180 3.545 4.050 3.885 ;
        RECT  3.820 3.545 4.050 4.250 ;
        RECT  5.150 3.625 5.490 4.250 ;
        RECT  3.820 4.020 5.490 4.250 ;
        RECT  2.430 0.980 2.770 1.320 ;
        RECT  5.150 0.980 5.490 1.320 ;
        RECT  0.805 1.090 5.490 1.320 ;
        RECT  0.805 1.090 1.035 1.840 ;
        RECT  0.660 1.500 1.035 1.840 ;
        RECT  3.995 1.090 4.225 2.630 ;
        RECT  3.995 2.400 4.660 2.630 ;
        RECT  4.430 2.400 4.660 3.790 ;
        RECT  4.430 3.505 4.770 3.790 ;
        RECT  0.805 1.090 4.80 1.320 ;
    END
END AO222X1

MACRO AO222X0
    CLASS CORE ;
    FOREIGN AO222X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.470 0.520 4.175 ;
        RECT  0.115 1.110 0.520 1.450 ;
        RECT  0.115 1.110 0.345 4.175 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.470 3.620 4.170 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.910 1.480 2.400 2.020 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.215 2.210 1.775 2.630 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.570 2.190 3.045 2.670 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.810 1.640 4.295 2.250 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.480 4.915 2.055 ;
        END
    END F
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  1.160 3.830 1.500 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.290 -0.400 3.630 0.790 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.780 2.850 1.120 3.190 ;
        RECT  0.780 2.960 2.410 3.190 ;
        RECT  2.180 2.960 2.410 4.250 ;
        RECT  2.180 3.930 3.030 4.250 ;
        RECT  2.780 2.900 3.120 3.240 ;
        RECT  2.780 3.010 4.080 3.240 ;
        RECT  3.850 3.010 4.080 4.250 ;
        RECT  3.850 3.930 4.360 4.250 ;
        RECT  2.040 0.910 2.380 1.250 ;
        RECT  4.520 0.910 4.860 1.250 ;
        RECT  0.755 1.020 4.860 1.250 ;
        RECT  0.755 1.020 0.985 2.270 ;
        RECT  0.575 1.930 0.985 2.270 ;
        RECT  3.350 1.020 3.580 2.780 ;
        RECT  3.350 2.550 4.595 2.780 ;
        RECT  4.310 2.550 4.595 3.130 ;
        RECT  0.755 1.020 3.40 1.250 ;
    END
END AO222X0

MACRO AO221X4
    CLASS CORE ;
    FOREIGN AO221X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 2.075 4.245 2.725 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.010 0.510 1.640 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.640 1.525 2.240 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 1.640 2.395 2.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.035 1.640 3.655 2.320 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 0.890 7.435 3.895 ;
        RECT  5.600 2.050 7.435 2.280 ;
        RECT  5.600 0.890 5.940 3.895 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.700 ;
        RECT  4.935 -0.400 5.220 1.700 ;
        RECT  3.325 -0.400 3.665 0.840 ;
        RECT  0.940 -0.400 1.280 1.410 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 2.640 6.660 5.280 ;
        RECT  4.935 2.640 5.220 5.280 ;
        RECT  1.675 3.610 2.015 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.905 3.150 2.775 3.380 ;
        RECT  0.905 3.150 1.245 4.180 ;
        RECT  2.435 3.150 2.775 4.180 ;
        RECT  0.180 2.690 3.610 2.920 ;
        RECT  0.180 2.690 0.520 4.180 ;
        RECT  3.270 2.690 3.610 4.180 ;
        RECT  2.135 1.070 4.705 1.410 ;
        RECT  4.475 1.945 5.370 2.285 ;
        RECT  4.475 1.070 4.705 3.185 ;
        RECT  4.075 2.955 4.705 3.185 ;
        RECT  4.075 2.955 4.415 4.180 ;
        RECT  0.180 2.690 2.40 2.920 ;
        RECT  2.135 1.070 3.30 1.410 ;
    END
END AO221X4

MACRO AO221X2
    CLASS CORE ;
    FOREIGN AO221X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.323  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.835 2.005 4.250 2.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.322  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.010 0.510 1.640 ;
        END
    END D
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.322  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.640 1.525 2.220 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.322  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 1.640 2.395 2.220 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.230 2.250 6.805 2.630 ;
        RECT  6.230 0.890 6.570 4.180 ;
        RECT  5.095 1.945 6.570 2.285 ;
        RECT  5.095 0.890 5.325 3.550 ;
        RECT  4.790 3.320 5.130 4.180 ;
        RECT  4.790 0.890 5.325 1.230 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.322  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.015 3.295 2.355 ;
        RECT  2.625 1.640 3.045 2.355 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.555 -0.400 5.850 1.230 ;
        RECT  3.325 -0.400 3.665 0.770 ;
        RECT  0.940 -0.400 1.280 1.340 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.510 3.840 5.850 5.280 ;
        RECT  5.555 3.260 5.850 5.280 ;
        RECT  1.675 3.610 2.015 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.905 3.150 2.775 3.380 ;
        RECT  0.905 3.150 1.245 4.180 ;
        RECT  2.435 3.150 2.775 4.180 ;
        RECT  0.180 2.690 3.610 2.920 ;
        RECT  0.180 2.690 0.520 4.180 ;
        RECT  3.270 2.690 3.610 4.180 ;
        RECT  2.135 1.000 4.425 1.340 ;
        RECT  4.195 1.000 4.425 1.775 ;
        RECT  4.195 1.545 4.865 1.775 ;
        RECT  4.480 1.545 4.865 1.885 ;
        RECT  4.480 1.545 4.710 3.090 ;
        RECT  4.035 2.860 4.710 3.090 ;
        RECT  4.035 2.860 4.375 4.180 ;
        RECT  0.180 2.690 2.20 2.920 ;
        RECT  2.135 1.000 3.50 1.340 ;
    END
END AO221X2

MACRO AO221X1
    CLASS CORE ;
    FOREIGN AO221X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.940 0.575 1.280 ;
        RECT  0.125 3.260 0.520 4.180 ;
        RECT  0.125 0.940 0.410 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.820 2.630 ;
        RECT  3.420 2.140 3.820 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.890 2.415 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.370 1.640 1.780 2.245 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.205 2.030 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.510 1.640 4.925 2.170 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  0.900 2.860 2.040 3.200 ;
        RECT  0.900 2.860 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.760 -0.400 4.100 0.950 ;
        RECT  1.055 -0.400 1.395 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.420 2.860 4.080 3.200 ;
        RECT  2.420 2.860 2.650 4.060 ;
        RECT  1.660 3.720 2.650 4.060 ;
        RECT  3.180 3.640 4.140 3.980 ;
        RECT  2.430 1.070 2.770 1.410 ;
        RECT  4.520 1.070 4.860 1.410 ;
        RECT  0.805 1.180 4.860 1.410 ;
        RECT  0.805 1.180 1.035 1.930 ;
        RECT  0.660 1.590 1.035 1.930 ;
        RECT  4.050 1.180 4.280 2.630 ;
        RECT  4.050 2.400 4.750 2.630 ;
        RECT  4.520 2.400 4.750 4.060 ;
        RECT  4.520 3.720 4.860 4.060 ;
        RECT  0.805 1.180 3.00 1.410 ;
    END
END AO221X1

MACRO AO221X0
    CLASS CORE ;
    FOREIGN AO221X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.930 0.520 4.250 ;
        RECT  0.125 1.030 0.520 1.495 ;
        RECT  0.125 1.030 0.355 4.250 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.117  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 1.640 2.395 2.525 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.117  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.315 1.640 1.775 2.225 ;
        END
    END A
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.117  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.030 3.035 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.117  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.640 3.675 2.375 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.117  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.400 4.285 2.120 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.290 3.930 1.630 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.090 -0.400 3.430 0.710 ;
        RECT  0.780 -0.400 1.120 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.045 2.860 3.965 3.200 ;
        RECT  2.320 2.860 2.660 3.790 ;
        RECT  2.060 0.830 2.400 1.170 ;
        RECT  3.890 0.680 4.230 1.170 ;
        RECT  0.755 0.940 4.230 1.170 ;
        RECT  0.755 0.940 0.985 2.115 ;
        RECT  0.585 1.775 0.815 3.660 ;
        RECT  0.585 3.430 2.090 3.660 ;
        RECT  1.860 3.430 2.090 4.250 ;
        RECT  3.890 3.930 4.230 4.250 ;
        RECT  1.860 4.020 4.230 4.250 ;
        RECT  1.045 2.860 2.40 3.200 ;
        RECT  0.755 0.940 3.80 1.170 ;
        RECT  1.860 4.020 3.40 4.250 ;
    END
END AO221X0

MACRO AO21X4
    CLASS CORE ;
    FOREIGN AO21X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.277  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.590 0.950 1.980 1.290 ;
        RECT  1.385 2.860 1.900 3.305 ;
        RECT  1.590 0.950 1.820 3.305 ;
        RECT  0.180 2.220 1.820 2.450 ;
        RECT  0.180 0.950 0.520 3.355 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 1.640 5.050 2.130 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.115 3.790 2.455 ;
        RECT  3.275 1.000 3.655 2.455 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.560 3.045 2.170 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  3.725 3.605 4.070 5.280 ;
        RECT  2.245 3.695 2.590 5.280 ;
        RECT  0.870 3.665 1.210 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.710 -0.400 5.050 1.410 ;
        RECT  2.485 -0.400 2.825 1.330 ;
        RECT  0.920 -0.400 1.260 1.290 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.970 3.145 4.770 3.375 ;
        RECT  4.430 3.145 4.770 4.155 ;
        RECT  2.970 3.145 3.310 4.175 ;
        RECT  3.910 0.950 4.250 1.290 ;
        RECT  2.050 2.035 2.390 2.385 ;
        RECT  2.160 2.035 2.390 2.915 ;
        RECT  4.020 0.950 4.250 2.915 ;
        RECT  2.160 2.685 5.490 2.915 ;
        RECT  5.145 2.685 5.490 4.180 ;
        RECT  2.160 2.685 4.90 2.915 ;
    END
END AO21X4

MACRO AO21X2
    CLASS CORE ;
    FOREIGN AO21X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.900 1.000 1.350 1.340 ;
        RECT  0.755 3.470 1.240 4.180 ;
        RECT  0.900 3.260 1.240 4.180 ;
        RECT  0.900 1.000 1.130 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 1.640 4.285 2.400 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.060 3.100 2.400 ;
        RECT  2.645 1.030 3.025 2.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.490 2.415 2.170 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  3.095 3.605 3.440 5.280 ;
        RECT  1.615 3.260 1.960 5.280 ;
        RECT  0.180 3.260 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  4.080 -0.400 4.420 1.390 ;
        RECT  1.855 -0.400 2.195 1.260 ;
        RECT  0.290 -0.400 0.630 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.340 3.145 4.140 3.375 ;
        RECT  2.340 3.145 2.680 4.175 ;
        RECT  3.800 3.145 4.140 4.180 ;
        RECT  3.280 0.965 3.620 1.305 ;
        RECT  1.420 2.540 1.760 2.915 ;
        RECT  3.390 0.965 3.620 2.915 ;
        RECT  1.420 2.685 4.860 2.915 ;
        RECT  4.515 2.685 4.860 4.190 ;
        RECT  1.420 2.685 3.40 2.915 ;
    END
END AO21X2

MACRO AO21X1
    CLASS CORE ;
    FOREIGN AO21X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.823  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.860 0.520 3.670 ;
        RECT  0.115 0.870 0.520 1.410 ;
        RECT  0.115 0.870 0.345 3.670 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 1.425 3.660 2.025 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 1.440 2.430 2.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.260 1.410 1.765 2.020 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  2.135 3.770 2.480 5.280 ;
        RECT  0.740 4.095 1.085 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.120 -0.400 3.460 1.180 ;
        RECT  0.980 -0.400 1.320 1.180 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.440 2.895 3.025 3.260 ;
        RECT  1.440 2.895 1.780 4.150 ;
        RECT  2.320 0.870 2.890 1.210 ;
        RECT  2.660 0.870 2.890 2.600 ;
        RECT  0.585 2.250 2.890 2.600 ;
        RECT  0.585 2.270 3.600 2.600 ;
        RECT  3.255 2.270 3.600 4.150 ;
        RECT  0.585 2.250 1.90 2.600 ;
        RECT  0.585 2.270 2.30 2.600 ;
    END
END AO21X1

MACRO AO21X0
    CLASS CORE ;
    FOREIGN AO21X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.582  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.930 0.520 4.250 ;
        RECT  0.115 0.630 0.520 1.410 ;
        RECT  0.115 0.630 0.345 4.250 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.295 2.160 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 1.030 3.025 1.865 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.121  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.535 0.630 1.970 0.880 ;
        RECT  1.385 1.030 1.765 1.410 ;
        RECT  1.535 0.630 1.765 1.410 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.980 3.965 1.790 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.560 -0.400 2.900 0.710 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.835 2.825 2.575 3.165 ;
        RECT  1.995 1.110 2.300 2.335 ;
        RECT  1.995 2.105 3.035 2.335 ;
        RECT  0.655 3.395 0.995 3.735 ;
        RECT  2.805 2.105 3.035 3.735 ;
        RECT  0.655 3.505 3.035 3.735 ;
        RECT  2.320 3.505 2.665 4.245 ;
        RECT  0.655 3.505 2.20 3.735 ;
    END
END AO21X0

MACRO AO211X4
    CLASS CORE ;
    FOREIGN AO211X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.190 2.630 ;
        RECT  1.850 2.175 2.190 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.545 2.630 ;
        RECT  0.115 1.915 0.525 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.470 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 0.890 6.120 3.895 ;
        RECT  4.340 2.250 6.120 2.630 ;
        RECT  4.340 0.890 4.680 3.895 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.450  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.420 2.175 2.975 2.660 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.060 2.860 5.400 5.280 ;
        RECT  3.665 2.640 3.960 5.280 ;
        RECT  0.940 3.350 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.060 -0.400 5.400 1.700 ;
        RECT  3.675 -0.400 3.960 1.700 ;
        RECT  3.620 -0.400 3.960 1.230 ;
        RECT  2.160 -0.400 2.445 1.320 ;
        RECT  0.180 -0.400 0.520 1.490 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.860 2.000 3.120 ;
        RECT  1.660 2.860 2.000 4.140 ;
        RECT  0.180 2.860 0.520 4.165 ;
        RECT  1.370 0.980 1.930 1.320 ;
        RECT  1.700 0.980 1.930 1.945 ;
        RECT  2.825 0.980 3.165 1.945 ;
        RECT  1.700 1.715 3.445 1.945 ;
        RECT  3.205 1.945 4.110 2.285 ;
        RECT  3.205 1.715 3.435 3.175 ;
        RECT  2.825 2.890 3.435 3.175 ;
        RECT  2.825 2.890 3.165 4.160 ;
    END
END AO211X4

MACRO AO211X2
    CLASS CORE ;
    FOREIGN AO211X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.190 2.630 ;
        RECT  1.850 2.120 2.190 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.010 0.525 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.470 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.899  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.245 2.250 4.920 2.630 ;
        RECT  4.245 1.010 4.585 4.175 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.420 2.120 3.035 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.965 3.255 5.305 5.280 ;
        RECT  3.525 3.320 3.865 5.280 ;
        RECT  0.940 3.320 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.965 -0.400 5.305 1.350 ;
        RECT  3.525 -0.400 3.865 1.350 ;
        RECT  2.160 -0.400 2.445 1.400 ;
        RECT  0.180 -0.400 0.520 1.490 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.860 2.000 3.090 ;
        RECT  0.180 2.860 0.520 3.760 ;
        RECT  1.660 2.860 2.000 3.760 ;
        RECT  1.370 1.060 1.930 1.400 ;
        RECT  1.700 1.060 1.930 1.880 ;
        RECT  2.825 1.060 3.165 1.880 ;
        RECT  1.700 1.650 4.015 1.880 ;
        RECT  3.265 1.650 4.015 1.990 ;
        RECT  3.265 1.650 3.495 3.090 ;
        RECT  2.825 2.860 3.495 3.090 ;
        RECT  2.825 2.860 3.165 3.760 ;
        RECT  1.700 1.650 3.80 1.880 ;
    END
END AO211X2

MACRO AO211X1
    CLASS CORE ;
    FOREIGN AO211X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.797  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.840 0.520 4.180 ;
        RECT  0.125 0.700 0.520 1.410 ;
        RECT  0.125 0.700 0.355 4.180 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.220  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.690 2.395 2.635 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.220  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.945 2.080 3.655 2.420 ;
        RECT  3.255 1.640 3.655 2.420 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.220  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.285 2.370 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.220  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.325 1.640 1.765 2.260 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  0.940 3.785 2.290 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.130 -0.400 3.470 0.710 ;
        RECT  0.940 -0.400 1.280 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.390 2.640 1.730 3.095 ;
        RECT  2.710 2.755 3.050 3.095 ;
        RECT  1.390 2.865 3.050 3.095 ;
        RECT  0.770 0.940 4.230 1.280 ;
        RECT  0.770 0.940 1.000 3.555 ;
        RECT  0.660 2.725 1.000 3.555 ;
        RECT  3.865 2.830 4.205 3.555 ;
        RECT  0.660 3.325 4.205 3.555 ;
        RECT  0.770 0.940 3.60 1.280 ;
        RECT  0.660 3.325 3.30 3.555 ;
    END
END AO211X1

MACRO AO211X0
    CLASS CORE ;
    FOREIGN AO211X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.670  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 3.965 0.520 4.250 ;
        RECT  0.125 0.630 0.520 1.410 ;
        RECT  0.125 0.630 0.355 4.250 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.975 1.995 2.395 2.635 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.215 1.640 1.745 2.260 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.640 3.025 2.420 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.112  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.820 3.655 2.630 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.290 3.965 1.630 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.560 -0.400 2.900 0.765 ;
        RECT  0.880 -0.400 1.220 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.045 2.850 1.360 3.190 ;
        RECT  1.045 2.960 2.660 3.190 ;
        RECT  2.320 2.960 2.660 3.790 ;
        RECT  3.260 0.630 3.600 1.355 ;
        RECT  0.755 1.015 3.600 1.355 ;
        RECT  0.755 1.015 0.985 2.070 ;
        RECT  0.585 1.840 0.815 3.735 ;
        RECT  0.585 3.395 0.940 3.735 ;
        RECT  0.585 3.505 2.090 3.735 ;
        RECT  1.860 3.505 2.090 4.250 ;
        RECT  3.060 3.930 3.400 4.250 ;
        RECT  1.860 4.020 3.400 4.250 ;
        RECT  0.755 1.015 2.20 1.355 ;
    END
END AO211X0

MACRO ANTENNACELLN5
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELLN5 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 0.970 0.590 1.470 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        END
    END vdd!
END ANTENNACELLN5

MACRO ANTENNACELLN25
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELLN25 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 0.970 0.590 1.470 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        END
    END vdd!
END ANTENNACELLN25

MACRO ANTENNACELLN2
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELLN2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 0.970 0.590 1.470 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        END
    END gnd!
END ANTENNACELLN2

MACRO ANTENNACELLN10
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELLN10 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 0.970 0.590 1.470 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        END
    END vdd!
END ANTENNACELLN10

MACRO ANTENNACELL5
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELL5 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.800 0.590 3.300 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        END
    END vdd!
END ANTENNACELL5

MACRO ANTENNACELL25
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELL25 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.750 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.800 0.590 3.300 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 15.750 0.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 15.750 5.280 ;
        END
    END vdd!
END ANTENNACELL25

MACRO ANTENNACELL2
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELL2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.800 0.590 3.300 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 1.260 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 1.260 0.400 ;
        END
    END gnd!
END ANTENNACELL2

MACRO ANTENNACELL10
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNACELL10 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNADIFFAREA 0.210  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.800 0.590 3.300 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        END
    END vdd!
END ANTENNACELL10

MACRO AND8X1
    CLASS CORE ;
    FOREIGN AND8X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.185 6.880 2.655 ;
        END
    END H
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.190 1.750 7.665 2.630 ;
        RECT  7.055 1.620 7.445 1.995 ;
        END
    END G
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.110 3.470 8.695 3.980 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.065 6.195 2.650 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.730 2.160 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.405 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.095 0.605 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.530  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.995 0.885 4.955 1.115 ;
        RECT  4.615 0.630 4.955 1.115 ;
        RECT  2.995 2.725 3.655 3.240 ;
        RECT  2.995 0.775 3.345 1.115 ;
        RECT  2.995 2.725 3.340 4.180 ;
        RECT  2.995 0.775 3.260 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 1.960 5.545 2.630 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  6.375 -0.400 6.715 1.690 ;
        RECT  3.805 -0.400 4.145 0.655 ;
        RECT  2.090 -0.400 2.430 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.540 3.640 7.880 5.280 ;
        RECT  6.160 2.900 6.500 5.280 ;
        RECT  4.575 3.360 4.915 5.280 ;
        RECT  2.250 2.995 2.590 5.280 ;
        RECT  0.770 3.735 1.110 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.370 0.520 1.820 ;
        RECT  2.425 1.480 2.765 1.820 ;
        RECT  0.180 1.590 2.765 1.820 ;
        RECT  0.935 1.590 1.165 3.310 ;
        RECT  0.180 2.970 1.870 3.310 ;
        RECT  5.145 1.330 5.485 1.670 ;
        RECT  4.685 1.345 5.485 1.670 ;
        RECT  3.665 1.690 4.915 2.030 ;
        RECT  4.685 1.345 4.915 3.130 ;
        RECT  4.685 2.900 5.750 3.130 ;
        RECT  5.410 2.900 5.750 3.240 ;
        RECT  8.120 0.630 8.655 0.970 ;
        RECT  8.120 0.630 8.460 3.240 ;
        RECT  6.880 2.900 8.640 3.240 ;
        RECT  0.180 1.590 1.50 1.820 ;
    END
END AND8X1

MACRO AND8X0
    CLASS CORE ;
    FOREIGN AND8X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.720 1.640 7.060 2.535 ;
        RECT  6.425 1.640 7.060 2.020 ;
        END
    END G
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 1.640 6.195 2.175 ;
        END
    END H
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.585 3.360 8.075 3.860 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.683  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.795 0.885 4.640 1.115 ;
        RECT  4.300 0.630 4.640 1.115 ;
        RECT  2.690 0.630 3.030 0.970 ;
        RECT  2.645 2.860 3.025 3.240 ;
        RECT  2.795 0.630 3.025 3.240 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.460 1.955 4.915 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.150 2.245 5.555 2.710 ;
        RECT  5.150 2.095 5.545 2.710 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.730 2.125 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.250 1.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.100 0.605 2.580 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.870 3.455 7.210 5.280 ;
        RECT  5.580 3.455 5.920 5.280 ;
        RECT  4.100 3.635 4.440 5.280 ;
        RECT  2.180 3.625 2.520 5.280 ;
        RECT  0.780 3.455 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  5.530 -0.400 6.350 1.410 ;
        RECT  3.490 -0.400 3.830 0.655 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.870 ;
        RECT  2.160 1.375 2.500 1.870 ;
        RECT  0.290 1.640 2.500 1.870 ;
        RECT  0.935 1.640 1.165 3.095 ;
        RECT  0.180 2.810 1.165 3.095 ;
        RECT  0.180 2.860 1.820 3.095 ;
        RECT  1.480 2.860 1.820 3.635 ;
        RECT  3.270 1.360 4.640 1.700 ;
        RECT  4.000 1.360 4.230 3.405 ;
        RECT  4.000 3.175 5.220 3.405 ;
        RECT  4.880 3.175 5.220 3.635 ;
        RECT  7.670 0.630 8.025 3.105 ;
        RECT  6.180 2.765 8.025 3.105 ;
        RECT  0.290 1.640 1.00 1.870 ;
    END
END AND8X0

MACRO AND7X1
    CLASS CORE ;
    FOREIGN AND7X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.095 0.605 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.390 0.915 ;
        RECT  0.755 0.630 1.135 1.360 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.730 2.160 2.395 2.630 ;
        END
    END C
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.220 6.905 2.655 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 1.960 5.545 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.065 6.195 2.650 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.530  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.960 0.885 4.955 1.115 ;
        RECT  4.615 0.630 4.955 1.115 ;
        RECT  2.995 2.685 3.655 3.240 ;
        RECT  2.995 2.685 3.340 4.180 ;
        RECT  2.995 0.800 3.300 4.180 ;
        RECT  2.960 0.800 3.300 1.140 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.190 1.750 7.610 2.270 ;
        RECT  7.055 1.620 7.445 1.995 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.375 -0.400 6.715 1.690 ;
        RECT  3.805 -0.400 4.145 0.655 ;
        RECT  2.045 -0.400 2.385 1.150 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.620 3.640 7.960 5.280 ;
        RECT  6.300 2.900 6.640 5.280 ;
        RECT  4.575 3.360 4.915 5.280 ;
        RECT  2.295 2.995 2.635 5.280 ;
        RECT  0.770 3.735 1.110 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.370 0.520 1.820 ;
        RECT  2.425 1.480 2.765 1.820 ;
        RECT  0.180 1.590 2.765 1.820 ;
        RECT  0.935 1.590 1.165 3.310 ;
        RECT  0.180 2.970 1.870 3.310 ;
        RECT  5.145 1.330 5.485 1.670 ;
        RECT  4.685 1.345 5.485 1.670 ;
        RECT  3.605 1.690 4.915 2.030 ;
        RECT  4.685 1.345 4.915 3.130 ;
        RECT  4.685 2.900 5.890 3.130 ;
        RECT  5.550 2.900 5.890 3.240 ;
        RECT  7.670 0.630 8.070 1.510 ;
        RECT  7.840 0.630 8.070 3.185 ;
        RECT  7.060 2.845 8.070 3.185 ;
        RECT  0.180 1.590 1.40 1.820 ;
    END
END AND7X1

MACRO AND7X0
    CLASS CORE ;
    FOREIGN AND7X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.100 0.605 2.580 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.220 1.410 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.730 2.100 2.395 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.150 2.075 5.565 2.675 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 1.620 6.865 2.220 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.120 6.195 2.630 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.079  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 1.960 4.915 2.660 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.683  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.690 0.885 4.640 1.115 ;
        RECT  4.300 0.630 4.640 1.115 ;
        RECT  2.690 0.630 3.030 1.115 ;
        RECT  2.645 2.820 3.025 3.240 ;
        RECT  2.690 0.630 2.920 3.240 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  5.590 -0.400 5.930 1.510 ;
        RECT  3.490 -0.400 3.830 0.655 ;
        RECT  1.640 -0.400 1.980 0.970 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.030 3.395 7.370 5.280 ;
        RECT  5.680 3.295 6.020 5.280 ;
        RECT  4.130 3.635 4.470 5.280 ;
        RECT  2.180 3.625 2.520 5.280 ;
        RECT  0.780 3.395 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.970 ;
        RECT  0.290 0.630 0.520 1.870 ;
        RECT  2.160 1.380 2.460 1.870 ;
        RECT  0.290 1.640 2.460 1.870 ;
        RECT  0.935 1.640 1.165 3.095 ;
        RECT  0.180 2.810 1.165 3.095 ;
        RECT  0.180 2.865 1.820 3.095 ;
        RECT  1.480 2.865 1.820 3.635 ;
        RECT  3.350 1.345 4.640 1.670 ;
        RECT  4.055 1.345 4.285 3.405 ;
        RECT  4.055 3.175 5.320 3.405 ;
        RECT  4.980 3.175 5.320 3.635 ;
        RECT  7.040 0.630 7.380 1.465 ;
        RECT  7.095 0.630 7.380 3.095 ;
        RECT  6.430 2.755 7.380 3.095 ;
        RECT  0.290 1.640 1.60 1.870 ;
    END
END AND7X0

MACRO AND6X4
    CLASS CORE ;
    FOREIGN AND6X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.180 0.655 2.710 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.250 5.325 2.660 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.285 2.365 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.905 1.640 5.545 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  9.545 1.130 9.955 4.105 ;
        RECT  8.280 2.365 9.955 2.615 ;
        RECT  8.120 2.850 8.510 4.105 ;
        RECT  8.280 1.130 8.510 4.105 ;
        RECT  8.120 1.130 8.510 1.470 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.150 2.415 2.745 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.345 2.180 1.765 2.790 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 10.080 5.280 ;
        RECT  8.840 2.850 9.180 5.280 ;
        RECT  7.360 4.170 7.700 5.280 ;
        RECT  6.040 3.825 6.380 5.280 ;
        RECT  4.795 3.825 5.135 5.280 ;
        RECT  2.130 3.820 2.470 5.280 ;
        RECT  0.970 3.815 1.310 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 10.080 0.400 ;
        RECT  8.840 -0.400 9.180 1.470 ;
        RECT  7.360 -0.400 7.700 0.710 ;
        RECT  6.180 -0.400 6.520 0.710 ;
        RECT  3.545 -0.400 3.885 1.250 ;
        RECT  1.840 -0.400 2.180 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.380 1.350 0.720 1.820 ;
        RECT  0.380 1.480 2.700 1.820 ;
        RECT  0.885 1.480 1.115 3.380 ;
        RECT  0.210 3.040 1.870 3.380 ;
        RECT  5.305 1.125 5.795 1.410 ;
        RECT  5.455 0.630 5.795 1.410 ;
        RECT  4.035 2.850 4.375 3.135 ;
        RECT  5.775 1.170 6.005 3.135 ;
        RECT  4.035 2.890 6.005 3.135 ;
        RECT  2.645 0.845 3.160 1.185 ;
        RECT  2.930 0.845 3.160 2.905 ;
        RECT  2.930 2.675 3.660 2.905 ;
        RECT  6.270 1.900 6.555 3.595 ;
        RECT  3.320 3.365 6.555 3.595 ;
        RECT  3.320 2.675 3.660 4.000 ;
        RECT  6.800 1.900 8.050 2.240 ;
        RECT  6.800 1.240 7.140 3.770 ;
        RECT  0.380 1.480 1.50 1.820 ;
        RECT  3.320 3.365 5.10 3.595 ;
    END
END AND6X4

MACRO AND6X2
    CLASS CORE ;
    FOREIGN AND6X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.975 0.505 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 3.470 2.030 4.220 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.115 2.120 5.565 2.640 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.528  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 4.515 1.870 ;
        RECT  4.170 1.130 4.515 1.870 ;
        RECT  3.410 1.640 3.750 3.790 ;
        RECT  3.275 1.640 3.750 2.020 ;
        RECT  2.645 0.790 2.985 1.870 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.620 6.175 2.830 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.353  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.925 3.470 7.435 4.250 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.280 3.525 6.620 5.280 ;
        RECT  4.560 2.860 4.900 5.280 ;
        RECT  2.260 2.860 2.600 5.280 ;
        RECT  0.740 4.095 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  4.890 -0.400 5.230 1.455 ;
        RECT  3.410 -0.400 3.750 1.270 ;
        RECT  1.840 -0.400 2.180 1.055 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.700 0.520 1.570 ;
        RECT  0.180 1.285 1.930 1.570 ;
        RECT  1.700 2.260 3.060 2.600 ;
        RECT  4.100 2.290 4.660 2.630 ;
        RECT  1.700 1.285 1.930 3.200 ;
        RECT  0.180 2.860 1.930 3.200 ;
        RECT  2.830 2.260 3.060 4.250 ;
        RECT  4.100 2.290 4.330 4.250 ;
        RECT  2.830 4.020 4.330 4.250 ;
        RECT  7.040 0.630 7.395 1.515 ;
        RECT  6.505 1.175 7.395 1.515 ;
        RECT  6.550 2.900 7.395 3.240 ;
        RECT  7.165 0.630 7.395 3.240 ;
        RECT  5.520 3.060 6.770 3.290 ;
        RECT  5.520 3.060 5.865 3.930 ;
    END
END AND6X2

MACRO AND6X1
    CLASS CORE ;
    FOREIGN AND6X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.845 2.300 5.545 2.640 ;
        RECT  5.165 1.640 5.545 2.640 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.650 2.205 2.395 2.630 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.245 0.950 ;
        RECT  0.755 0.630 1.135 1.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.175 0.630 2.655 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.872  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.860 3.025 3.960 ;
        RECT  2.730 0.820 2.960 3.960 ;
        RECT  2.560 0.820 2.960 1.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.960 4.515 2.630 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.775 2.045 6.185 2.640 ;
        END
    END F
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 1.690 ;
        RECT  3.280 -0.400 3.620 1.120 ;
        RECT  1.840 -0.400 2.180 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.020 3.640 5.360 5.280 ;
        RECT  3.820 3.640 4.160 5.280 ;
        RECT  1.300 3.735 1.640 5.280 ;
        RECT  0.180 3.735 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.630 0.520 0.960 ;
        RECT  0.290 0.630 0.520 1.870 ;
        RECT  2.160 1.480 2.500 1.870 ;
        RECT  0.290 1.640 2.500 1.870 ;
        RECT  0.935 1.640 1.165 3.295 ;
        RECT  0.740 2.955 2.400 3.295 ;
        RECT  3.440 1.350 4.540 1.690 ;
        RECT  3.190 1.690 3.670 2.030 ;
        RECT  3.440 1.350 3.670 3.210 ;
        RECT  3.440 2.870 6.120 3.210 ;
        RECT  0.290 1.640 1.40 1.870 ;
        RECT  3.440 2.870 5.60 3.210 ;
    END
END AND6X1

MACRO AND6X0
    CLASS CORE ;
    FOREIGN AND6X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.150 1.625 5.550 2.245 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.598  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.210 2.860 3.655 3.535 ;
        RECT  3.210 1.170 3.440 3.535 ;
        RECT  2.870 1.170 3.440 1.510 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.245 0.505 2.875 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.420 0.915 ;
        RECT  0.755 0.630 1.135 1.410 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.100 1.990 2.630 ;
        END
    END F
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.890 2.090 4.305 2.660 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.575 5.015 3.340 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.125 4.225 5.465 5.280 ;
        RECT  3.725 4.225 4.065 5.280 ;
        RECT  2.180 4.010 2.520 5.280 ;
        RECT  0.780 3.890 1.120 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  3.740 -0.400 4.080 1.510 ;
        RECT  2.020 -0.400 2.360 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.520 1.870 ;
        RECT  0.180 1.640 0.965 1.870 ;
        RECT  0.735 1.640 0.965 3.590 ;
        RECT  0.180 3.250 0.965 3.590 ;
        RECT  2.330 1.890 2.670 3.535 ;
        RECT  0.180 3.305 2.670 3.535 ;
        RECT  0.180 3.305 1.820 3.590 ;
        RECT  1.480 3.305 1.820 4.130 ;
        RECT  5.485 1.025 6.065 1.365 ;
        RECT  5.725 3.280 6.065 3.995 ;
        RECT  5.780 1.025 6.065 3.995 ;
        RECT  2.930 3.765 6.065 3.995 ;
        RECT  2.930 3.765 3.270 4.130 ;
        RECT  4.425 3.765 4.765 4.160 ;
        RECT  0.180 3.305 1.40 3.535 ;
        RECT  2.930 3.765 5.80 3.995 ;
    END
END AND6X0

MACRO AND5X4
    CLASS CORE ;
    FOREIGN AND5X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.450 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.345 2.180 1.765 2.790 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.250 4.285 2.900 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.180 0.655 2.710 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.275 1.640 4.915 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.915 1.130 9.325 4.105 ;
        RECT  7.650 2.365 9.325 2.615 ;
        RECT  7.475 2.850 7.880 4.105 ;
        RECT  7.650 1.130 7.880 4.105 ;
        RECT  7.490 1.130 7.880 1.470 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.150 2.415 2.745 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 9.450 5.280 ;
        RECT  8.210 2.850 8.550 5.280 ;
        RECT  6.730 4.170 7.070 5.280 ;
        RECT  5.410 3.825 5.750 5.280 ;
        RECT  4.035 3.825 4.375 5.280 ;
        RECT  2.130 3.820 2.470 5.280 ;
        RECT  0.970 3.815 1.310 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 9.450 0.400 ;
        RECT  8.210 -0.400 8.550 1.470 ;
        RECT  6.730 -0.400 7.070 0.710 ;
        RECT  5.550 -0.400 5.890 0.710 ;
        RECT  3.445 -0.400 3.785 1.650 ;
        RECT  1.840 -0.400 2.180 0.950 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.380 1.350 0.720 1.820 ;
        RECT  0.380 1.480 2.700 1.820 ;
        RECT  0.885 1.480 1.115 3.380 ;
        RECT  0.210 3.040 1.870 3.380 ;
        RECT  4.675 1.125 5.165 1.410 ;
        RECT  4.825 0.630 5.165 1.410 ;
        RECT  5.145 1.170 5.375 3.135 ;
        RECT  4.595 2.850 5.375 3.135 ;
        RECT  2.645 0.815 3.160 1.155 ;
        RECT  2.930 0.815 3.160 2.905 ;
        RECT  2.930 2.675 3.660 2.905 ;
        RECT  5.605 1.900 5.890 3.595 ;
        RECT  3.320 3.365 5.890 3.595 ;
        RECT  3.320 2.675 3.660 4.000 ;
        RECT  6.155 1.900 7.420 2.240 ;
        RECT  6.155 1.225 6.510 3.770 ;
        RECT  0.380 1.480 1.40 1.820 ;
        RECT  3.320 3.365 4.40 3.595 ;
    END
END AND5X4

MACRO AND5X2
    CLASS CORE ;
    FOREIGN AND5X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.900 6.270 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.110 1.640 5.545 2.550 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.470 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 3.470 2.150 4.220 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.530 0.525 2.125 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.469  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.835 1.640 4.475 1.870 ;
        RECT  4.135 1.100 4.475 1.870 ;
        RECT  3.530 1.640 3.870 3.790 ;
        RECT  3.275 1.640 3.870 2.020 ;
        RECT  2.835 0.810 3.065 1.870 ;
        RECT  2.560 0.810 3.065 1.150 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.855 -0.400 5.195 1.410 ;
        RECT  3.375 -0.400 3.715 1.320 ;
        RECT  1.800 -0.400 2.140 1.230 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.540 6.750 5.280 ;
        RECT  4.680 2.780 5.020 5.280 ;
        RECT  2.380 2.780 2.720 5.280 ;
        RECT  0.900 3.320 1.205 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.960 0.985 1.300 ;
        RECT  0.755 0.960 0.985 1.710 ;
        RECT  0.755 1.480 2.605 1.710 ;
        RECT  1.920 1.480 2.605 1.820 ;
        RECT  1.920 2.250 3.300 2.480 ;
        RECT  4.100 2.210 4.780 2.550 ;
        RECT  0.180 2.860 2.150 3.090 ;
        RECT  1.920 1.480 2.150 3.200 ;
        RECT  1.620 2.860 2.150 3.200 ;
        RECT  0.180 2.860 0.520 3.700 ;
        RECT  3.070 2.250 3.300 4.250 ;
        RECT  4.100 2.210 4.330 4.250 ;
        RECT  3.070 4.020 4.330 4.250 ;
        RECT  6.425 0.630 6.765 1.545 ;
        RECT  5.995 1.205 6.765 1.545 ;
        RECT  6.500 0.630 6.765 3.230 ;
        RECT  5.690 3.000 6.765 3.230 ;
        RECT  5.690 3.000 6.045 3.920 ;
    END
END AND5X2

MACRO AND5X1
    CLASS CORE ;
    FOREIGN AND5X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.920 3.690 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.145 2.045 5.555 2.640 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.200 2.250 1.765 2.735 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.130 0.510 2.745 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.028  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.165 0.820 2.485 1.160 ;
        RECT  2.000 2.640 2.395 3.960 ;
        RECT  2.165 0.820 2.395 3.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.215 2.300 4.915 2.640 ;
        RECT  4.535 1.640 4.915 2.640 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.150 -0.400 5.490 1.690 ;
        RECT  2.865 -0.400 3.205 1.120 ;
        RECT  1.275 -0.400 1.615 1.160 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.390 3.640 4.730 5.280 ;
        RECT  3.190 3.640 3.530 5.280 ;
        RECT  1.300 3.735 1.640 5.280 ;
        RECT  0.180 3.735 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.640 0.520 0.980 ;
        RECT  0.290 0.640 0.520 1.800 ;
        RECT  1.595 1.460 1.935 1.800 ;
        RECT  0.290 1.570 1.935 1.800 ;
        RECT  0.740 1.570 0.970 3.295 ;
        RECT  0.740 2.955 1.080 3.295 ;
        RECT  2.815 1.350 3.910 1.690 ;
        RECT  2.670 1.690 3.045 2.030 ;
        RECT  2.815 1.350 3.045 3.210 ;
        RECT  2.815 2.870 5.490 3.210 ;
        RECT  2.815 2.870 4.30 3.210 ;
    END
END AND5X1

MACRO AND5X0
    CLASS CORE ;
    FOREIGN AND5X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.830 2.250 2.395 2.685 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.195 1.640 1.780 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.245 0.505 2.875 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.566  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.210 2.860 3.655 3.535 ;
        RECT  3.210 1.160 3.440 3.535 ;
        RECT  3.050 1.160 3.440 1.500 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.760 5.015 3.240 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.170 4.305 2.705 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.920 -0.400 4.260 1.500 ;
        RECT  2.180 -0.400 2.520 1.500 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.125 4.225 5.465 5.280 ;
        RECT  3.725 4.225 4.065 5.280 ;
        RECT  2.180 4.110 2.520 5.280 ;
        RECT  0.780 3.900 1.120 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.360 0.965 1.700 ;
        RECT  2.625 2.240 2.965 2.590 ;
        RECT  0.735 1.360 0.965 3.590 ;
        RECT  0.180 3.250 0.965 3.590 ;
        RECT  2.625 2.240 2.855 3.535 ;
        RECT  0.180 3.305 2.855 3.535 ;
        RECT  0.180 3.305 1.820 3.590 ;
        RECT  1.480 3.305 1.820 4.240 ;
        RECT  5.150 1.160 5.490 1.500 ;
        RECT  5.245 1.160 5.490 3.995 ;
        RECT  2.930 3.765 5.490 3.995 ;
        RECT  4.425 3.765 4.765 4.230 ;
        RECT  2.930 3.765 3.270 4.250 ;
        RECT  0.180 3.305 1.20 3.535 ;
        RECT  2.930 3.765 4.80 3.995 ;
    END
END AND5X0

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.820 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.130 1.415 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.655 2.900 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.180 0.520 2.790 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.645 1.640 4.285 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  8.285 1.130 8.695 4.105 ;
        RECT  7.060 2.365 8.695 2.615 ;
        RECT  6.845 2.850 7.290 4.105 ;
        RECT  7.060 1.130 7.290 4.105 ;
        RECT  6.860 1.130 7.290 1.470 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.820 5.280 ;
        RECT  7.580 2.850 7.920 5.280 ;
        RECT  6.100 4.170 6.440 5.280 ;
        RECT  4.780 3.825 5.120 5.280 ;
        RECT  3.405 3.825 3.745 5.280 ;
        RECT  1.500 3.820 1.840 5.280 ;
        RECT  0.180 3.080 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.820 0.400 ;
        RECT  7.580 -0.400 7.920 1.470 ;
        RECT  6.100 -0.400 6.440 0.710 ;
        RECT  4.920 -0.400 5.260 0.710 ;
        RECT  2.815 -0.400 3.155 1.650 ;
        RECT  1.210 -0.400 1.550 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.350 0.520 1.825 ;
        RECT  0.180 1.540 2.070 1.825 ;
        RECT  1.645 1.540 2.070 1.880 ;
        RECT  1.645 1.540 1.875 3.380 ;
        RECT  0.900 3.040 1.875 3.380 ;
        RECT  4.045 1.125 4.535 1.410 ;
        RECT  4.195 0.630 4.535 1.410 ;
        RECT  4.515 1.170 4.745 3.135 ;
        RECT  3.965 2.850 4.745 3.135 ;
        RECT  2.015 0.815 2.585 1.155 ;
        RECT  2.355 0.815 2.585 3.010 ;
        RECT  2.355 2.675 3.030 3.010 ;
        RECT  4.975 1.900 5.260 3.595 ;
        RECT  2.690 3.365 5.260 3.595 ;
        RECT  2.690 2.675 3.030 4.000 ;
        RECT  5.525 1.900 6.830 2.240 ;
        RECT  5.525 1.225 5.880 3.770 ;
        RECT  2.690 3.365 4.80 3.595 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.250 1.470 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.480 2.125 4.915 2.630 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.575 0.525 2.175 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.700 5.725 2.270 ;
        RECT  5.165 1.640 5.595 2.270 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.525  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.310 3.870 1.650 ;
        RECT  2.770 1.310 3.115 3.790 ;
        RECT  2.645 1.310 3.115 2.020 ;
        RECT  2.050 1.310 3.870 1.560 ;
        RECT  2.050 0.815 2.390 1.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 2.960 6.120 5.280 ;
        RECT  3.960 2.775 4.300 5.280 ;
        RECT  1.620 3.540 1.960 5.280 ;
        RECT  0.180 3.075 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.250 -0.400 4.590 1.520 ;
        RECT  2.770 -0.400 3.110 1.080 ;
        RECT  1.330 -0.400 1.670 1.155 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 0.880 1.030 1.220 ;
        RECT  0.800 0.880 1.030 2.020 ;
        RECT  0.800 1.790 2.150 2.020 ;
        RECT  1.810 1.790 2.150 2.130 ;
        RECT  3.500 2.160 4.070 2.500 ;
        RECT  1.810 1.790 2.040 3.310 ;
        RECT  0.900 3.080 2.540 3.310 ;
        RECT  0.900 3.080 1.240 4.000 ;
        RECT  2.310 3.080 2.540 4.250 ;
        RECT  3.500 2.160 3.730 4.250 ;
        RECT  2.310 4.020 3.730 4.250 ;
        RECT  5.780 0.630 6.185 1.470 ;
        RECT  5.955 0.630 6.185 2.730 ;
        RECT  5.145 2.500 6.185 2.730 ;
        RECT  5.145 2.500 5.375 3.745 ;
        RECT  5.035 2.860 5.375 3.745 ;
    END
END AND4X2

MACRO AND4X1
    CLASS CORE ;
    FOREIGN AND4X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.525 2.870 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.115 1.470 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 2.250 3.675 2.920 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.102  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.490 2.640 3.025 3.960 ;
        RECT  2.490 1.045 2.720 3.960 ;
        RECT  2.380 1.045 2.720 1.385 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.250 4.335 2.850 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.495 4.170 4.835 5.280 ;
        RECT  3.295 4.170 3.635 5.280 ;
        RECT  1.390 3.890 1.730 5.280 ;
        RECT  0.180 3.890 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.195 -0.400 3.535 1.385 ;
        RECT  1.480 -0.400 1.820 1.385 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.165 0.520 1.885 ;
        RECT  0.180 1.655 2.260 1.885 ;
        RECT  1.700 1.655 2.260 2.030 ;
        RECT  1.700 1.655 1.930 3.450 ;
        RECT  0.790 3.110 1.930 3.450 ;
        RECT  4.425 1.165 4.795 2.020 ;
        RECT  2.950 1.690 4.795 2.020 ;
        RECT  4.565 1.165 4.795 3.680 ;
        RECT  3.895 3.340 4.795 3.680 ;
        RECT  0.180 1.655 1.80 1.885 ;
    END
END AND4X1

MACRO AND4X0
    CLASS CORE ;
    FOREIGN AND4X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.541  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.580 2.860 3.025 3.535 ;
        RECT  2.580 1.170 2.810 3.535 ;
        RECT  2.395 1.170 2.810 1.510 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.250 0.525 2.870 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.200 1.415 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.275 1.905 3.675 2.645 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.090 4.330 2.740 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  4.495 4.225 4.835 5.280 ;
        RECT  3.095 4.225 3.435 5.280 ;
        RECT  1.590 4.170 1.930 5.280 ;
        RECT  0.180 3.885 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.195 -0.400 3.535 1.510 ;
        RECT  1.480 -0.400 1.820 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 1.170 0.520 1.970 ;
        RECT  0.180 1.740 1.875 1.970 ;
        RECT  1.645 2.215 2.260 2.550 ;
        RECT  1.645 1.740 1.875 3.590 ;
        RECT  0.790 3.250 1.875 3.590 ;
        RECT  4.425 1.170 4.790 1.510 ;
        RECT  3.895 3.515 4.235 3.995 ;
        RECT  4.560 1.170 4.790 3.995 ;
        RECT  2.340 3.765 4.790 3.995 ;
        RECT  2.340 3.765 2.680 4.220 ;
        RECT  2.340 3.765 3.30 3.995 ;
    END
END AND4X0

MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.170 0.580 2.525 ;
        RECT  0.115 2.170 0.510 2.710 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 2.860 6.805 3.955 ;
        RECT  6.410 0.905 6.750 3.955 ;
        RECT  4.970 2.085 6.750 2.365 ;
        RECT  4.970 0.905 5.310 3.955 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 1.640 2.395 2.315 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.702  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.090 0.630 3.430 2.520 ;
        RECT  1.330 0.630 3.430 0.860 ;
        RECT  1.220 1.640 1.560 2.520 ;
        RECT  1.330 0.630 1.560 2.520 ;
        RECT  0.755 1.640 1.560 2.020 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 2.700 6.030 5.280 ;
        RECT  4.180 4.170 4.520 5.280 ;
        RECT  2.900 3.210 3.240 5.280 ;
        RECT  1.460 3.210 1.800 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.245 ;
        RECT  3.940 -0.400 4.280 1.505 ;
        RECT  0.270 -0.400 0.610 1.305 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.180 1.090 2.855 1.410 ;
        RECT  2.625 1.090 2.855 2.980 ;
        RECT  4.425 1.685 4.740 2.980 ;
        RECT  0.740 2.750 4.740 2.980 ;
        RECT  0.740 2.750 1.080 3.620 ;
        RECT  2.180 2.750 2.520 3.620 ;
        RECT  3.620 2.750 3.960 3.620 ;
        RECT  0.740 2.750 3.70 2.980 ;
    END
END AND3X4

MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.953  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.240 3.870 ;
        RECT  0.755 0.860 1.240 1.200 ;
        RECT  0.755 0.860 0.995 3.870 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.850 2.170 4.295 2.720 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.635 2.115 3.070 2.675 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.351  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 1.640 2.405 2.350 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  3.100 3.410 3.440 5.280 ;
        RECT  1.620 3.410 1.960 5.280 ;
        RECT  0.180 2.930 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  1.770 -0.400 2.110 1.165 ;
        RECT  0.180 -0.400 0.520 1.210 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  3.390 0.700 3.730 1.570 ;
        RECT  1.225 2.260 1.565 3.180 ;
        RECT  3.390 0.700 3.620 3.180 ;
        RECT  1.225 2.950 4.200 3.180 ;
        RECT  2.340 2.950 2.680 3.870 ;
        RECT  3.860 2.950 4.200 3.870 ;
        RECT  1.225 2.950 3.30 3.180 ;
    END
END AND3X2

MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.061  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.910 0.520 4.250 ;
        RECT  0.115 0.820 0.520 1.410 ;
        RECT  0.115 0.820 0.345 4.250 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.655 1.510 3.035 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.680 2.860 2.395 3.240 ;
        RECT  1.680 2.090 1.965 3.240 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.140 1.460 1.765 1.800 ;
        RECT  1.415 1.030 1.765 1.800 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.980 4.170 2.320 5.280 ;
        RECT  0.880 4.170 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  0.900 -0.400 1.185 1.160 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.195 0.820 2.820 1.160 ;
        RECT  2.195 0.820 2.425 2.630 ;
        RECT  0.580 2.090 0.920 2.430 ;
        RECT  2.195 2.400 2.855 2.630 ;
        RECT  0.690 2.090 0.920 3.700 ;
        RECT  2.625 2.400 2.855 3.700 ;
        RECT  0.690 3.470 2.970 3.700 ;
        RECT  1.430 3.470 1.770 3.930 ;
        RECT  2.630 3.470 2.970 3.960 ;
        RECT  0.690 3.470 1.70 3.700 ;
    END
END AND3X1

MACRO AND3X0
    CLASS CORE ;
    FOREIGN AND3X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.750 2.115 1.145 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 1.955 2.850 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.005 3.030 2.635 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.487  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.930 0.600 4.250 ;
        RECT  0.115 1.170 0.520 2.020 ;
        RECT  0.115 1.170 0.355 4.250 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.930 3.810 2.270 5.280 ;
        RECT  0.830 3.070 1.070 5.280 ;
        RECT  0.585 3.070 1.070 3.410 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.010 -0.400 1.350 0.900 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.185 1.170 2.810 1.510 ;
        RECT  2.185 1.170 2.415 3.500 ;
        RECT  1.300 3.160 2.415 3.500 ;
        RECT  1.300 3.270 2.860 3.500 ;
        RECT  2.630 3.270 2.860 4.150 ;
        RECT  2.630 3.810 2.970 4.150 ;
        RECT  1.300 3.160 1.640 4.190 ;
    END
END AND3X0

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.100 1.740 2.630 2.080 ;
        RECT  2.100 0.710 2.330 2.080 ;
        RECT  0.750 0.710 2.330 0.940 ;
        RECT  0.115 1.630 0.980 1.860 ;
        RECT  0.750 0.710 0.980 1.860 ;
        RECT  0.115 1.630 0.560 2.030 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.648  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.175 1.305 2.695 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.249  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.020 2.250 5.550 2.630 ;
        RECT  5.020 2.250 5.360 4.100 ;
        RECT  4.760 0.900 5.100 2.480 ;
        RECT  3.580 2.250 5.550 2.480 ;
        RECT  3.580 2.250 3.920 4.100 ;
        RECT  3.580 0.900 3.810 4.100 ;
        RECT  3.320 0.900 3.810 1.240 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  4.295 2.850 4.650 5.280 ;
        RECT  2.820 2.850 3.160 5.280 ;
        RECT  1.300 4.170 1.640 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.040 -0.400 4.380 1.240 ;
        RECT  2.560 -0.400 2.900 1.510 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.370 1.170 1.765 1.510 ;
        RECT  3.010 2.280 3.350 2.620 ;
        RECT  1.535 2.335 3.350 2.620 ;
        RECT  1.535 1.170 1.765 3.475 ;
        RECT  0.740 3.135 2.400 3.475 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.000 2.200 2.535 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.324  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.900 2.150 3.655 2.490 ;
        RECT  3.275 1.640 3.655 2.490 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.470 1.240 4.010 ;
        RECT  0.835 3.090 1.240 4.010 ;
        RECT  0.835 1.040 1.240 1.380 ;
        RECT  0.835 1.040 1.065 4.010 ;
        END
    END Q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  1.660 -0.400 2.000 1.410 ;
        RECT  0.180 -0.400 0.520 1.380 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  3.140 3.090 3.480 5.280 ;
        RECT  1.660 3.350 2.000 5.280 ;
        RECT  0.180 3.090 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.815 0.995 3.190 1.335 ;
        RECT  2.815 0.995 3.045 1.920 ;
        RECT  1.380 1.690 3.045 1.920 ;
        RECT  1.380 1.690 1.740 2.030 ;
        RECT  1.510 1.690 1.740 3.120 ;
        RECT  1.510 2.890 2.760 3.120 ;
        RECT  2.420 2.890 2.760 4.010 ;
    END
END AND2X2

MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.059  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.905 0.520 4.245 ;
        RECT  0.115 1.030 0.520 1.530 ;
        RECT  0.115 1.030 0.345 4.245 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.210 1.640 1.765 2.460 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.238  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.995 2.120 2.395 3.240 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  2.000 4.170 2.340 5.280 ;
        RECT  0.880 4.170 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.875 -0.400 1.215 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.750 1.180 2.340 1.410 ;
        RECT  2.000 1.180 2.340 1.520 ;
        RECT  0.575 2.120 0.980 2.460 ;
        RECT  0.750 1.180 0.980 3.820 ;
        RECT  0.750 3.590 1.790 3.820 ;
        RECT  1.450 3.590 1.790 3.930 ;
    END
END AND2X1

MACRO AND2X0
    CLASS CORE ;
    FOREIGN AND2X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.190 2.245 1.770 2.665 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.104  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 2.120 2.395 3.240 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.723  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 3.470 0.520 4.180 ;
        RECT  0.115 0.630 0.520 0.970 ;
        RECT  0.115 0.630 0.345 4.180 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  1.730 3.890 2.070 5.280 ;
        RECT  0.880 3.890 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  0.970 -0.400 1.310 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  2.000 1.170 2.340 1.510 ;
        RECT  0.575 1.280 2.340 1.510 ;
        RECT  0.575 1.280 0.860 3.220 ;
        RECT  0.575 2.990 1.780 3.220 ;
        RECT  1.480 2.990 1.780 3.430 ;
    END
END AND2X0

MACRO AN33X4
    CLASS CORE ;
    FOREIGN AN33X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.390 0.525 3.245 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.205 2.470 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.421  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.910 1.560 2.510 2.020 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.325 2.250 3.780 2.710 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.040  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.880 2.920 7.380 3.260 ;
        RECT  5.595 1.485 7.375 1.715 ;
        RECT  7.035 0.890 7.375 1.715 ;
        RECT  6.425 1.485 6.805 3.260 ;
        RECT  5.595 0.890 5.935 1.715 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.585 2.250 3.095 2.710 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 2.250 2.055 2.710 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.460 3.560 6.800 5.280 ;
        RECT  5.225 3.555 5.565 5.280 ;
        RECT  1.325 3.680 1.675 5.280 ;
        RECT  0.175 3.680 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.315 -0.400 6.655 1.230 ;
        RECT  4.930 -0.400 5.215 1.230 ;
        RECT  3.565 -0.400 3.905 0.835 ;
        RECT  0.235 -0.400 0.580 1.470 ;
        RECT  0.235 -0.400 0.525 1.520 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.755 2.940 3.615 3.280 ;
        RECT  1.890 0.955 3.345 1.295 ;
        RECT  3.115 0.955 3.345 1.970 ;
        RECT  3.115 1.720 4.240 1.970 ;
        RECT  4.010 2.120 4.525 2.460 ;
        RECT  4.010 1.720 4.240 4.020 ;
        RECT  2.605 3.680 4.240 4.020 ;
        RECT  4.155 1.150 4.700 1.490 ;
        RECT  4.470 1.460 4.985 1.690 ;
        RECT  4.755 1.945 6.075 2.285 ;
        RECT  4.755 1.460 4.985 3.260 ;
        RECT  4.590 2.915 4.985 3.260 ;
        RECT  0.755 2.940 2.10 3.280 ;
    END
END AN33X4

MACRO AN33X2
    CLASS CORE ;
    FOREIGN AN33X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.390 0.505 3.245 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.610 1.575 2.020 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.640 2.740 2.020 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.210 1.620 3.810 2.020 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.250 3.320 2.720 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.335 2.250 2.055 2.720 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.750 6.190 3.560 ;
        RECT  5.960 1.250 6.190 3.560 ;
        RECT  5.850 1.250 6.190 1.590 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.960 6.750 5.280 ;
        RECT  5.090 3.960 5.430 5.280 ;
        RECT  1.300 3.890 1.640 5.280 ;
        RECT  0.175 3.890 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 0.720 ;
        RECT  5.285 -0.400 5.630 0.725 ;
        RECT  3.780 -0.400 4.120 0.910 ;
        RECT  0.235 -0.400 0.580 1.020 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.950 3.600 3.290 ;
        RECT  2.000 2.950 2.340 4.230 ;
        RECT  2.160 0.700 2.500 1.390 ;
        RECT  2.160 1.140 4.285 1.390 ;
        RECT  4.040 1.945 4.455 2.285 ;
        RECT  4.040 1.140 4.285 4.230 ;
        RECT  2.695 3.890 4.285 4.230 ;
        RECT  4.530 1.250 4.915 1.590 ;
        RECT  4.685 1.945 5.730 2.285 ;
        RECT  4.685 1.250 4.915 3.560 ;
        RECT  4.530 2.750 4.915 3.560 ;
        RECT  0.740 2.950 2.30 3.290 ;
        RECT  2.160 1.140 3.20 1.390 ;
    END
END AN33X2

MACRO AN33X1
    CLASS CORE ;
    FOREIGN AN33X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.390 0.540 3.245 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.445 1.575 2.020 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.640 2.740 2.020 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.495 1.640 3.825 2.040 ;
        RECT  3.090 1.640 3.825 2.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.836  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.605 3.680 4.285 4.020 ;
        RECT  4.055 1.030 4.285 4.020 ;
        RECT  2.160 1.030 4.285 1.410 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.250 3.320 2.720 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.335 2.250 2.055 2.720 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.325 3.680 1.675 5.280 ;
        RECT  0.175 3.680 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.780 -0.400 4.120 0.710 ;
        RECT  0.235 -0.400 0.580 1.280 ;
        RECT  0.235 -0.400 0.525 1.520 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.770 2.950 3.615 3.290 ;
        RECT  0.770 2.950 2.80 3.290 ;
    END
END AN33X1

MACRO AN33X0
    CLASS CORE ;
    FOREIGN AN33X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.045 0.525 2.635 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.540 1.315 2.005 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.510 2.555 2.010 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.090 1.555 3.665 2.020 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.134  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.695 3.530 4.285 3.920 ;
        RECT  4.055 1.030 4.285 3.920 ;
        RECT  3.905 1.030 4.285 1.410 ;
        RECT  1.935 1.030 4.285 1.280 ;
        RECT  1.935 0.680 2.275 1.280 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.250 3.235 2.580 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.355 2.240 2.045 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.295 3.580 1.645 5.280 ;
        RECT  0.175 3.580 0.525 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.605 -0.400 3.945 0.800 ;
        RECT  0.265 -0.400 0.610 1.020 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.735 2.790 1.075 3.130 ;
        RECT  3.260 2.810 3.600 3.130 ;
        RECT  0.735 2.860 3.600 3.130 ;
        RECT  1.995 2.860 2.335 3.920 ;
        RECT  0.735 2.860 2.60 3.130 ;
    END
END AN33X0

MACRO AN333X1
    CLASS CORE ;
    FOREIGN AN333X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 1.640 4.285 2.200 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 1.640 3.035 2.125 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.135 1.030 1.765 1.410 ;
        RECT  1.135 1.030 1.475 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.850 2.245 2.395 2.630 ;
        RECT  1.850 2.120 2.250 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 1.955 3.655 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.666  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.400 2.860 6.815 4.180 ;
        RECT  6.585 1.030 6.815 4.180 ;
        RECT  2.315 1.180 6.815 1.410 ;
        RECT  6.220 1.030 6.815 1.410 ;
        RECT  5.020 2.860 6.815 3.200 ;
        RECT  2.315 1.070 2.655 1.410 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 1.640 6.320 2.115 ;
        END
    END G
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.515 1.965 4.935 2.630 ;
        END
    END J
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.760 5.565 2.630 ;
        END
    END H
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.120 0.760 2.630 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  4.215 -0.400 4.555 0.950 ;
        RECT  0.180 -0.400 0.520 1.510 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  1.620 3.370 1.960 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 4.020 3.140 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  2.340 2.860 4.020 3.200 ;
        RECT  3.010 3.680 6.030 4.020 ;
        RECT  0.900 2.860 3.60 3.140 ;
        RECT  3.010 3.680 5.90 4.020 ;
    END
END AN333X1

MACRO AN333X0
    CLASS CORE ;
    FOREIGN AN333X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.930 1.590 5.555 2.020 ;
        END
    END H
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.780 1.560 4.350 2.020 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 1.350 3.035 2.020 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.135 1.640 1.775 2.020 ;
        RECT  1.135 1.640 1.475 2.120 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.825 2.245 2.415 2.660 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.085 2.245 3.670 2.660 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.160 0.760 2.630 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.040  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.415 0.940 6.815 1.410 ;
        RECT  4.860 2.910 6.645 3.200 ;
        RECT  6.415 0.940 6.645 3.200 ;
        RECT  6.180 2.860 6.645 3.200 ;
        RECT  3.340 0.940 6.815 1.180 ;
        RECT  5.880 0.680 6.220 1.180 ;
        RECT  2.315 0.680 3.570 1.020 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.250 6.185 2.630 ;
        RECT  5.900 1.855 6.185 2.630 ;
        END
    END G
    PIN J
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.355 2.250 4.925 2.680 ;
        END
    END J
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  3.980 -0.400 4.320 0.710 ;
        RECT  0.655 -0.400 0.995 1.020 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  1.460 3.680 1.800 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  0.900 2.890 3.880 3.200 ;
        RECT  2.980 3.680 5.760 4.020 ;
        RECT  0.900 2.890 2.80 3.200 ;
        RECT  2.980 3.680 4.20 4.020 ;
    END
END AN333X0

MACRO AN332X1
    CLASS CORE ;
    FOREIGN AN332X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.935  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.055 2.830 6.185 3.060 ;
        RECT  5.955 1.030 6.185 3.060 ;
        RECT  2.315 1.070 6.185 1.410 ;
        RECT  5.590 1.030 6.185 1.410 ;
        RECT  5.055 2.830 5.400 3.610 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.120 0.760 2.630 ;
        END
    END A
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.465  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.760 4.935 2.630 ;
        END
    END G
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.446  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 1.640 5.690 2.115 ;
        END
    END H
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 1.640 4.285 2.160 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.580 1.640 3.035 2.105 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.135 1.030 1.765 1.410 ;
        RECT  1.135 1.030 1.475 2.120 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.850 2.245 2.395 2.630 ;
        RECT  1.850 2.120 2.350 2.630 ;
        END
    END C
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 2.010 3.655 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  1.620 3.320 1.960 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  4.215 -0.400 4.555 0.840 ;
        RECT  0.180 -0.400 0.520 1.580 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 4.020 3.090 ;
        RECT  0.900 2.860 1.240 3.200 ;
        RECT  2.340 2.860 4.020 3.200 ;
        RECT  3.010 3.840 6.120 4.180 ;
        RECT  0.900 2.860 3.80 3.090 ;
        RECT  3.010 3.840 5.30 4.180 ;
    END
END AN332X1

MACRO AN332X0
    CLASS CORE ;
    FOREIGN AN332X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.085 0.525 2.645 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.530 1.220 2.020 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.470 2.550 1.970 ;
        END
    END F
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.720 4.305 2.630 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.085 1.475 3.655 1.970 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.798  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.590 2.745 5.555 3.085 ;
        RECT  5.325 0.680 5.555 3.085 ;
        RECT  5.165 0.680 5.555 1.410 ;
        RECT  1.930 0.940 5.555 1.180 ;
        RECT  5.150 0.680 5.555 1.180 ;
        RECT  1.930 0.680 2.270 1.180 ;
        END
    END Q
    PIN H
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.095 2.140 ;
        END
    END H
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.200 3.270 2.580 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.375 2.200 2.010 2.580 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.700 -0.400 4.040 0.710 ;
        RECT  0.270 -0.400 0.610 1.020 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  1.300 3.565 1.640 5.280 ;
        RECT  0.180 3.565 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.810 3.600 3.150 ;
        RECT  2.000 2.810 2.340 3.905 ;
        RECT  2.700 3.565 5.490 3.905 ;
        RECT  0.740 2.810 2.70 3.150 ;
        RECT  2.700 3.565 4.30 3.905 ;
    END
END AN332X0

MACRO AN331X1
    CLASS CORE ;
    FOREIGN AN331X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 2.010 3.655 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.690  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.140 2.860 5.555 4.140 ;
        RECT  5.325 0.940 5.555 4.140 ;
        RECT  2.315 1.170 5.555 1.410 ;
        RECT  4.975 0.940 5.555 1.410 ;
        RECT  2.315 1.070 2.655 1.410 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.120 0.760 2.630 ;
        END
    END A
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.060 2.145 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 1.640 4.285 2.305 ;
        END
    END D
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.483  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.640 3.025 2.190 ;
        END
    END F
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.135 1.030 1.765 1.410 ;
        RECT  1.135 1.030 1.475 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.850 2.245 2.395 2.630 ;
        RECT  1.850 2.120 2.250 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  1.620 3.425 1.960 5.280 ;
        RECT  0.180 2.860 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  4.215 -0.400 4.555 0.940 ;
        RECT  0.180 -0.400 0.520 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 4.020 3.195 ;
        RECT  3.010 3.680 4.690 4.020 ;
        RECT  0.900 2.860 3.70 3.195 ;
    END
END AN331X1

MACRO AN331X0
    CLASS CORE ;
    FOREIGN AN331X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.040 0.525 2.635 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.525 1.235 2.020 ;
        END
    END B
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.410 2.550 1.970 ;
        END
    END F
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.090 1.470 3.660 1.970 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.918  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 3.565 4.915 3.905 ;
        RECT  4.685 0.680 4.915 3.905 ;
        RECT  4.535 0.680 4.915 1.410 ;
        RECT  1.930 0.940 4.915 1.180 ;
        RECT  4.400 0.680 4.915 1.180 ;
        RECT  1.930 0.680 2.270 1.180 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.144  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 2.250 4.455 2.630 ;
        RECT  4.120 1.765 4.455 2.630 ;
        END
    END G
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.640 2.200 3.270 2.580 ;
        RECT  2.640 2.200 3.210 2.585 ;
        END
    END E
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.200 2.010 2.585 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.600 -0.400 3.940 0.710 ;
        RECT  0.240 -0.400 0.580 1.020 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  1.300 3.565 1.640 5.280 ;
        RECT  0.180 3.565 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.815 3.600 3.155 ;
        RECT  2.000 2.815 2.340 3.905 ;
        RECT  2.700 3.565 4.160 3.905 ;
        RECT  0.740 2.815 2.90 3.155 ;
    END
END AN331X0

MACRO AN32X4
    CLASS CORE ;
    FOREIGN AN32X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.205 2.470 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.435 2.250 2.055 2.720 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.250 3.155 2.720 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.040  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.970 1.485 6.750 1.715 ;
        RECT  6.410 0.890 6.750 1.715 ;
        RECT  5.210 2.920 6.710 3.260 ;
        RECT  5.795 1.485 6.175 3.260 ;
        RECT  4.970 0.890 5.310 1.715 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.735 1.640 2.395 2.020 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.390 0.525 3.245 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.230 ;
        RECT  4.305 -0.400 4.590 1.230 ;
        RECT  2.990 -0.400 3.330 0.780 ;
        RECT  0.175 -0.400 0.520 1.525 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.790 3.560 6.130 5.280 ;
        RECT  4.555 3.555 4.895 5.280 ;
        RECT  1.325 3.680 1.675 5.280 ;
        RECT  0.180 3.680 0.525 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.755 2.950 2.245 3.290 ;
        RECT  1.955 2.950 2.245 4.020 ;
        RECT  1.955 3.680 3.560 4.020 ;
        RECT  1.760 0.970 2.855 1.310 ;
        RECT  2.625 0.970 2.855 2.020 ;
        RECT  2.625 1.790 3.615 2.020 ;
        RECT  3.385 2.120 3.845 2.460 ;
        RECT  3.385 1.790 3.615 3.250 ;
        RECT  2.630 2.950 3.615 3.250 ;
        RECT  3.530 1.105 4.070 1.445 ;
        RECT  3.840 1.105 4.070 1.690 ;
        RECT  3.840 1.460 4.305 1.690 ;
        RECT  4.075 1.945 5.235 2.285 ;
        RECT  4.075 1.460 4.305 3.260 ;
        RECT  3.920 2.915 4.305 3.260 ;
    END
END AN32X4

MACRO AN32X2
    CLASS CORE ;
    FOREIGN AN32X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.445 1.430 2.020 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.335 2.250 2.055 2.720 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.192  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.250 3.195 2.720 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.750 5.560 3.560 ;
        RECT  5.330 1.250 5.560 3.560 ;
        RECT  5.220 1.250 5.560 1.590 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.192  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 1.635 2.645 2.020 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.390 0.540 3.245 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 0.720 ;
        RECT  4.660 -0.400 5.000 0.720 ;
        RECT  3.255 -0.400 3.595 0.925 ;
        RECT  0.175 -0.400 0.520 1.050 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 3.960 6.120 5.280 ;
        RECT  4.460 3.960 4.800 5.280 ;
        RECT  1.335 2.950 1.685 5.280 ;
        RECT  0.175 4.170 0.525 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  2.040 0.700 2.385 1.405 ;
        RECT  2.040 1.155 3.655 1.405 ;
        RECT  3.425 1.945 3.865 2.285 ;
        RECT  3.425 1.155 3.655 3.545 ;
        RECT  2.660 3.205 3.655 3.545 ;
        RECT  3.900 1.360 4.325 1.700 ;
        RECT  4.095 1.945 5.100 2.285 ;
        RECT  4.095 1.360 4.325 2.980 ;
        RECT  3.900 2.640 4.325 2.980 ;
    END
END AN32X2

MACRO AN32X1
    CLASS CORE ;
    FOREIGN AN32X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.445 1.430 2.020 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.335 2.250 2.055 2.720 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.250 3.195 2.720 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.244  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.950 3.655 3.290 ;
        RECT  3.425 1.030 3.655 3.290 ;
        RECT  2.040 1.030 3.655 1.410 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.406  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.010 1.640 2.645 2.020 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.422  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.390 0.540 3.245 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.255 -0.400 3.595 0.800 ;
        RECT  0.175 -0.400 0.520 1.525 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.325 3.680 1.675 5.280 ;
        RECT  0.175 3.680 0.525 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.770 2.950 2.245 3.290 ;
        RECT  1.955 2.950 2.245 4.020 ;
        RECT  1.955 3.680 3.560 4.020 ;
    END
END AN32X1

MACRO AN32X0
    CLASS CORE ;
    FOREIGN AN32X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.110 0.525 2.665 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.585 1.320 2.020 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.158  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.350 2.475 2.020 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.535  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.660 2.860 3.655 3.160 ;
        RECT  3.425 1.030 3.655 3.160 ;
        RECT  3.275 1.030 3.655 1.410 ;
        RECT  2.705 1.030 3.655 1.270 ;
        RECT  2.705 0.735 2.935 1.270 ;
        RECT  1.930 0.735 2.935 1.020 ;
        RECT  1.930 0.680 2.270 1.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.158  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.560 2.250 3.195 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.020 2.640 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.300 3.590 1.640 5.280 ;
        RECT  0.180 3.590 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  3.165 -0.400 3.505 0.710 ;
        RECT  0.240 -0.400 0.580 1.020 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.820 1.080 3.160 ;
        RECT  0.740 2.870 2.330 3.160 ;
        RECT  2.100 2.870 2.330 3.930 ;
        RECT  2.100 3.590 3.560 3.930 ;
    END
END AN32X0

MACRO AN322X1
    CLASS CORE ;
    FOREIGN AN322X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.685 2.250 2.395 2.630 ;
        RECT  1.685 2.120 2.025 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 1.995 3.655 2.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.757  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.495 2.760 5.545 3.100 ;
        RECT  5.315 0.700 5.545 3.100 ;
        RECT  1.930 1.170 5.545 1.410 ;
        RECT  5.000 0.700 5.545 1.410 ;
        RECT  1.930 1.070 2.270 1.410 ;
        END
    END Q
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.305 2.200 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.355 1.640 3.025 2.020 ;
        END
    END E
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.995 1.640 1.335 2.460 ;
        RECT  0.755 1.640 1.335 2.020 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.050 0.525 2.635 ;
        END
    END A
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 1.640 5.085 2.200 ;
        END
    END G
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.300 -0.400 4.115 0.940 ;
        RECT  0.180 -0.400 0.520 1.580 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  1.330 3.580 1.670 5.280 ;
        RECT  0.180 3.580 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.755 2.860 3.430 3.200 ;
        RECT  2.515 3.580 5.485 3.920 ;
        RECT  0.755 2.860 2.70 3.200 ;
        RECT  2.515 3.580 4.80 3.920 ;
    END
END AN322X1

MACRO AN322X0
    CLASS CORE ;
    FOREIGN AN322X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.080 0.525 2.665 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.555 1.220 1.970 ;
        RECT  0.755 1.555 1.160 2.100 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.455 2.550 1.805 ;
        RECT  2.015 1.455 2.445 1.970 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.795 1.640 4.325 2.160 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.781  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.590 2.810 5.545 3.100 ;
        RECT  5.315 0.980 5.545 3.100 ;
        RECT  1.930 0.940 5.340 1.180 ;
        RECT  5.165 0.980 5.545 1.410 ;
        RECT  5.000 0.680 5.340 1.180 ;
        RECT  1.930 0.680 2.270 1.180 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.255 4.995 2.580 ;
        RECT  4.655 1.675 4.995 2.580 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.157  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.595 2.150 3.220 2.505 ;
        RECT  2.595 2.150 3.035 2.620 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.162  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.380 2.200 1.990 2.620 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  3.160 -0.400 3.990 0.710 ;
        RECT  0.270 -0.400 0.610 1.020 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  1.300 3.570 1.640 5.280 ;
        RECT  0.180 3.570 0.520 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.750 1.080 3.090 ;
        RECT  0.740 2.850 3.600 3.090 ;
        RECT  3.260 2.810 3.600 3.140 ;
        RECT  2.000 2.850 3.600 3.140 ;
        RECT  2.000 2.850 2.340 3.910 ;
        RECT  2.700 3.570 5.490 3.910 ;
        RECT  0.740 2.850 2.30 3.090 ;
        RECT  2.700 3.570 4.20 3.910 ;
    END
END AN322X0

MACRO AN321X4
    CLASS CORE ;
    FOREIGN AN321X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.050 0.525 2.635 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.995 1.640 1.335 2.500 ;
        RECT  0.755 1.640 1.335 2.020 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.355 1.640 3.025 2.020 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.365 2.170 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.952  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.510 2.920 8.010 3.260 ;
        RECT  6.400 1.360 8.010 1.700 ;
        RECT  7.055 1.360 7.435 3.260 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 1.995 3.655 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.685 2.250 2.395 2.630 ;
        RECT  1.685 2.120 2.025 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.090 3.560 7.430 5.280 ;
        RECT  5.855 3.555 6.195 5.280 ;
        RECT  1.330 3.580 1.670 5.280 ;
        RECT  0.180 3.580 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.035 -0.400 7.375 1.130 ;
        RECT  5.810 -0.400 6.150 1.080 ;
        RECT  3.500 -0.400 3.840 0.940 ;
        RECT  0.180 -0.400 0.520 1.580 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.755 2.860 3.430 3.200 ;
        RECT  2.515 3.580 4.130 3.920 ;
        RECT  1.930 1.070 2.270 1.410 ;
        RECT  4.505 0.700 4.860 1.410 ;
        RECT  1.930 1.170 4.860 1.410 ;
        RECT  4.630 2.120 4.990 2.460 ;
        RECT  4.630 0.700 4.860 3.100 ;
        RECT  4.520 2.760 4.860 3.100 ;
        RECT  5.220 1.945 6.500 2.285 ;
        RECT  5.220 1.360 5.560 3.260 ;
        RECT  0.755 2.860 2.80 3.200 ;
        RECT  1.930 1.170 3.60 1.410 ;
    END
END AN321X4

MACRO AN321X2
    CLASS CORE ;
    FOREIGN AN321X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.050 0.525 2.635 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.995 1.640 1.335 2.460 ;
        RECT  0.755 1.640 1.335 2.020 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.217  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.355 1.640 3.025 2.020 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.420 2.200 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.425 2.750 6.820 3.560 ;
        RECT  6.590 1.250 6.820 3.560 ;
        RECT  6.480 1.250 6.820 1.590 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.217  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 2.080 3.655 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.685 2.250 2.395 2.630 ;
        RECT  1.685 2.120 2.025 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  7.040 3.960 7.380 5.280 ;
        RECT  5.720 3.960 6.060 5.280 ;
        RECT  1.300 3.760 1.640 5.280 ;
        RECT  0.180 3.760 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  7.040 -0.400 7.380 0.720 ;
        RECT  5.920 -0.400 6.260 0.720 ;
        RECT  3.480 -0.400 3.820 0.940 ;
        RECT  0.180 -0.400 0.520 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.860 3.600 3.200 ;
        RECT  1.995 2.860 2.340 4.100 ;
        RECT  2.700 3.760 4.100 4.100 ;
        RECT  1.930 1.070 2.270 1.410 ;
        RECT  4.460 1.070 4.880 1.410 ;
        RECT  1.930 1.170 4.880 1.410 ;
        RECT  4.650 1.945 5.050 2.285 ;
        RECT  4.650 1.070 4.880 4.100 ;
        RECT  4.465 3.760 4.880 4.100 ;
        RECT  5.160 1.275 5.510 1.615 ;
        RECT  5.280 1.945 6.360 2.285 ;
        RECT  5.280 1.275 5.510 3.560 ;
        RECT  5.160 2.750 5.510 3.560 ;
        RECT  0.740 2.860 2.40 3.200 ;
        RECT  1.930 1.170 3.90 1.410 ;
    END
END AN321X2

MACRO AN321X1
    CLASS CORE ;
    FOREIGN AN321X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 2.160 0.545 2.635 ;
        RECT  0.120 2.120 0.540 2.635 ;
        RECT  0.120 2.050 0.525 2.635 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.995 1.640 1.335 2.500 ;
        RECT  0.755 1.640 1.335 2.020 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.355 1.640 3.025 2.020 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.428  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.905 1.640 4.365 2.200 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.720  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.520 2.760 4.915 3.100 ;
        RECT  4.685 0.700 4.915 3.100 ;
        RECT  1.930 1.170 4.915 1.410 ;
        RECT  4.505 0.700 4.915 1.410 ;
        RECT  1.930 1.070 2.270 1.410 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.466  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 1.995 3.655 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.482  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.685 2.250 2.395 2.630 ;
        RECT  1.685 2.120 2.025 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  1.330 3.580 1.670 5.280 ;
        RECT  0.180 3.580 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.500 -0.400 3.840 0.940 ;
        RECT  0.180 -0.400 0.520 1.580 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.755 2.860 3.430 3.200 ;
        RECT  2.515 3.580 4.130 3.920 ;
        RECT  0.755 2.860 2.40 3.200 ;
    END
END AN321X1

MACRO AN321X0
    CLASS CORE ;
    FOREIGN AN321X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.045 0.580 2.630 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 0.630 1.440 0.945 ;
        RECT  0.755 0.630 1.135 1.410 ;
        END
    END B
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.005 3.460 2.435 4.040 ;
        END
    END E
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.167  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.755 3.920 3.605 4.250 ;
        RECT  3.275 3.470 3.605 4.250 ;
        END
    END F
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.764  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.860 3.680 4.285 4.020 ;
        RECT  3.950 1.360 4.285 4.020 ;
        RECT  3.890 1.360 4.285 2.020 ;
        RECT  1.960 1.360 4.285 1.590 ;
        RECT  1.960 1.360 2.300 1.700 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.184  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.880 3.280 2.220 ;
        RECT  2.645 1.880 3.025 2.630 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.985 1.990 2.325 ;
        RECT  1.385 1.985 1.765 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.300 3.560 1.640 5.280 ;
        RECT  0.180 3.560 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.220 -0.400 3.560 1.025 ;
        RECT  0.180 -0.400 0.520 1.700 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.800 1.080 3.140 ;
        RECT  2.060 2.720 2.400 3.140 ;
        RECT  3.380 2.720 3.720 3.140 ;
        RECT  0.740 2.910 3.720 3.140 ;
        RECT  0.740 2.910 2.60 3.140 ;
    END
END AN321X0

MACRO AN31X4
    CLASS CORE ;
    FOREIGN AN31X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.105 0.525 2.830 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.360 1.470 2.700 ;
        RECT  0.755 1.640 1.155 2.700 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.210 0.890 6.550 3.560 ;
        RECT  4.880 2.250 6.550 2.630 ;
        RECT  4.770 2.750 5.110 3.560 ;
        RECT  4.880 0.890 5.110 3.560 ;
        RECT  4.770 0.890 5.110 1.700 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.520 1.900 2.045 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.625 2.760 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.490 2.860 5.830 5.280 ;
        RECT  4.050 2.750 4.390 5.280 ;
        RECT  1.470 3.800 1.810 5.280 ;
        RECT  0.180 3.800 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.490 -0.400 5.830 1.700 ;
        RECT  4.050 -0.400 4.390 1.700 ;
        RECT  2.630 -0.400 2.970 1.180 ;
        RECT  0.180 -0.400 0.520 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.890 2.990 2.390 3.330 ;
        RECT  1.795 0.940 2.360 1.280 ;
        RECT  2.130 0.940 2.360 1.645 ;
        RECT  2.130 1.415 3.085 1.645 ;
        RECT  2.855 1.945 3.255 2.285 ;
        RECT  2.855 1.415 3.085 4.180 ;
        RECT  2.630 3.840 3.085 4.180 ;
        RECT  3.330 0.890 3.715 1.700 ;
        RECT  3.485 1.945 4.650 2.285 ;
        RECT  3.485 0.890 3.715 3.920 ;
        RECT  3.330 2.640 3.715 3.920 ;
    END
END AN31X4

MACRO AN31X2
    CLASS CORE ;
    FOREIGN AN31X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.105 0.525 2.730 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.390 1.470 2.730 ;
        RECT  0.755 1.640 1.155 2.730 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.535 2.750 4.930 3.560 ;
        RECT  4.700 1.250 4.930 3.560 ;
        RECT  4.590 1.250 4.930 1.590 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.605 1.845 2.135 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.178  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.535 1.460 3.025 2.020 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 3.960 5.490 5.280 ;
        RECT  3.830 3.960 4.170 5.280 ;
        RECT  1.400 3.030 1.740 5.280 ;
        RECT  0.180 4.170 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.150 -0.400 5.490 0.720 ;
        RECT  4.030 -0.400 4.370 0.720 ;
        RECT  2.630 -0.400 2.970 0.950 ;
        RECT  0.180 -0.400 0.520 1.040 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  1.795 0.730 2.305 1.070 ;
        RECT  2.075 0.730 2.305 2.480 ;
        RECT  2.075 2.250 3.250 2.480 ;
        RECT  2.660 2.250 3.250 2.520 ;
        RECT  2.660 2.250 3.000 4.230 ;
        RECT  3.270 1.360 3.710 1.700 ;
        RECT  3.480 1.945 4.470 2.285 ;
        RECT  3.480 1.360 3.710 3.005 ;
        RECT  3.270 2.750 3.610 3.560 ;
    END
END AN31X2

MACRO AN31X1
    CLASS CORE ;
    FOREIGN AN31X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.105 0.525 2.730 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.360 1.470 2.700 ;
        RECT  0.755 1.640 1.155 2.700 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.971  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.525 2.970 4.180 ;
        RECT  2.075 2.525 2.970 2.755 ;
        RECT  1.795 0.940 2.395 1.410 ;
        RECT  2.075 0.940 2.305 2.755 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.420  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 1.640 1.845 2.130 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.378  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.535 1.640 3.025 2.180 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  1.470 3.800 1.810 5.280 ;
        RECT  0.180 3.800 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 1.280 ;
        RECT  0.180 -0.400 0.520 1.510 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.890 2.990 2.390 3.330 ;
    END
END AN31X1

MACRO AN31X0
    CLASS CORE ;
    FOREIGN AN31X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.105 0.525 2.670 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.155 2.430 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.667  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 2.410 2.970 2.980 ;
        RECT  2.075 2.410 2.970 2.640 ;
        RECT  2.015 1.030 2.395 1.600 ;
        RECT  2.075 1.030 2.305 2.640 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.146  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.640 3.025 2.180 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.166  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.120 1.845 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.460 3.900 1.555 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.220 -0.400 2.560 0.740 ;
        RECT  0.180 -0.400 0.520 1.480 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.475 2.910 2.300 3.150 ;
        RECT  0.475 2.910 0.815 3.250 ;
        RECT  2.070 2.910 2.300 3.770 ;
        RECT  2.070 3.430 2.410 3.770 ;
    END
END AN31X0

MACRO AN311X4
    CLASS CORE ;
    FOREIGN AN311X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.640 0.525 2.235 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.100 1.470 2.440 ;
        RECT  0.755 1.640 1.135 2.440 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.040 0.810 7.380 3.560 ;
        RECT  5.600 2.250 7.380 2.630 ;
        RECT  5.600 0.810 5.940 3.560 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 1.640 2.395 2.160 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.080 3.025 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 2.080 3.655 2.630 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 7.560 5.280 ;
        RECT  6.320 2.860 6.660 5.280 ;
        RECT  4.895 2.945 5.220 5.280 ;
        RECT  1.620 3.330 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 7.560 0.400 ;
        RECT  6.320 -0.400 6.660 1.620 ;
        RECT  4.895 -0.400 5.220 1.620 ;
        RECT  2.860 -0.400 3.200 0.840 ;
        RECT  0.180 -0.400 0.520 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 2.690 3.100 ;
        RECT  0.900 2.860 1.240 4.140 ;
        RECT  2.320 2.860 2.690 4.140 ;
        RECT  2.060 1.070 3.850 1.410 ;
        RECT  3.620 1.295 4.115 1.635 ;
        RECT  3.885 1.940 4.205 2.285 ;
        RECT  3.885 1.295 4.115 3.090 ;
        RECT  3.490 2.860 4.115 3.090 ;
        RECT  3.490 2.860 3.830 3.200 ;
        RECT  4.160 0.685 4.665 1.040 ;
        RECT  4.435 1.945 5.370 2.285 ;
        RECT  4.435 0.685 4.665 3.600 ;
        RECT  4.160 3.370 4.500 4.180 ;
    END
END AN311X4

MACRO AN311X2
    CLASS CORE ;
    FOREIGN AN311X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.560 0.525 2.230 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.430 2.230 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.225  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 2.170 2.395 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.985 3.025 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.255 1.985 3.615 2.630 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.690 2.860 6.175 3.560 ;
        RECT  5.690 1.250 6.030 3.560 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 2.750 6.750 5.280 ;
        RECT  4.970 2.750 5.310 5.280 ;
        RECT  1.620 3.330 1.960 5.280 ;
        RECT  0.180 3.140 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.410 -0.400 6.750 1.565 ;
        RECT  4.965 -0.400 5.310 1.565 ;
        RECT  2.570 -0.400 2.910 0.710 ;
        RECT  0.180 -0.400 0.520 1.290 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 2.690 3.100 ;
        RECT  0.900 2.860 1.240 3.505 ;
        RECT  2.320 2.860 2.690 3.505 ;
        RECT  1.760 0.940 4.075 1.280 ;
        RECT  3.845 1.945 4.205 2.285 ;
        RECT  3.845 0.940 4.075 3.500 ;
        RECT  3.490 3.160 4.075 3.500 ;
        RECT  4.305 1.255 4.665 1.595 ;
        RECT  4.435 1.945 5.460 2.285 ;
        RECT  4.435 1.255 4.665 3.560 ;
        RECT  4.305 2.750 4.665 3.560 ;
        RECT  1.760 0.940 3.50 1.280 ;
    END
END AN311X2

MACRO AN311X1
    CLASS CORE ;
    FOREIGN AN311X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.620 0.525 2.235 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.060 1.470 2.400 ;
        RECT  0.755 1.640 1.135 2.400 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.600  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.885 0.940 4.285 1.410 ;
        RECT  3.490 2.250 4.115 2.590 ;
        RECT  3.885 0.940 4.115 2.590 ;
        RECT  2.060 0.940 4.285 1.280 ;
        RECT  3.490 2.250 3.830 4.180 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.464  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.860 1.620 2.395 2.105 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 2.170 3.025 2.630 ;
        RECT  2.625 2.120 2.985 2.630 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.410  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.210 1.510 3.655 2.020 ;
        END
    END E
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.620 3.330 1.960 5.280 ;
        RECT  0.180 2.640 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  2.860 -0.400 3.200 0.710 ;
        RECT  0.180 -0.400 0.520 1.390 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 2.860 2.690 3.100 ;
        RECT  0.900 2.860 1.240 4.140 ;
        RECT  2.320 2.860 2.690 4.140 ;
    END
END AN311X1

MACRO AN311X0
    CLASS CORE ;
    FOREIGN AN311X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.500 0.555 2.055 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 3.320 1.295 3.850 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.178  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.675 2.480 2.580 ;
        END
    END D
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.178  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.020 3.325 3.655 3.850 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.819  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 2.690 3.655 3.030 ;
        RECT  3.425 1.005 3.655 3.030 ;
        RECT  1.860 1.005 3.655 1.360 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.202  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.260 1.600 1.785 2.020 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.570 3.660 1.910 5.280 ;
        RECT  0.180 3.660 0.520 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.660 -0.400 3.000 0.710 ;
        RECT  0.180 -0.400 0.520 0.715 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 2.720 1.080 3.060 ;
        RECT  0.740 2.820 2.610 3.060 ;
        RECT  2.270 2.820 2.610 4.000 ;
    END
END AN311X0

MACRO AN22X4
    CLASS CORE ;
    FOREIGN AN22X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.210 0.890 6.550 3.895 ;
        RECT  4.770 2.250 6.550 2.630 ;
        RECT  4.770 0.890 5.110 3.895 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.580 1.500 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.285 2.250 1.885 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.580 2.625 2.060 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.190 0.600 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.490 2.860 5.830 5.280 ;
        RECT  4.050 2.640 4.390 5.280 ;
        RECT  0.760 3.550 1.100 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.490 -0.400 5.830 1.700 ;
        RECT  4.050 -0.400 4.390 1.700 ;
        RECT  2.565 -0.400 2.905 0.780 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.900 1.675 3.240 ;
        RECT  1.335 2.900 1.675 3.880 ;
        RECT  1.335 3.540 2.985 3.880 ;
        RECT  1.370 1.010 3.085 1.350 ;
        RECT  2.855 1.945 3.255 2.285 ;
        RECT  2.855 1.010 3.085 3.235 ;
        RECT  2.055 2.895 3.085 3.235 ;
        RECT  3.330 0.780 3.715 1.700 ;
        RECT  3.485 1.945 4.540 2.285 ;
        RECT  3.485 0.780 3.715 4.180 ;
        RECT  3.330 2.640 3.715 4.180 ;
    END
END AN22X4

MACRO AN22X2
    CLASS CORE ;
    FOREIGN AN22X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.060 2.785 5.545 3.705 ;
        RECT  5.315 1.240 5.545 3.705 ;
        RECT  5.060 1.240 5.545 1.580 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.630 1.500 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.085 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.630 2.805 2.020 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.190 0.600 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 2.785 6.120 5.280 ;
        RECT  4.340 2.785 4.680 5.280 ;
        RECT  0.745 3.820 1.085 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 1.580 ;
        RECT  4.340 -0.400 4.680 1.580 ;
        RECT  2.645 -0.400 2.985 0.830 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.910 1.845 3.250 ;
        RECT  1.505 2.910 1.845 4.160 ;
        RECT  1.505 3.820 3.260 4.160 ;
        RECT  1.410 1.060 3.350 1.400 ;
        RECT  3.120 2.090 3.500 2.430 ;
        RECT  3.120 1.060 3.350 3.250 ;
        RECT  2.225 2.910 3.350 3.250 ;
        RECT  3.580 1.240 3.960 1.580 ;
        RECT  3.730 2.090 5.085 2.430 ;
        RECT  3.730 1.240 3.960 3.705 ;
        RECT  3.620 2.785 3.960 3.705 ;
    END
END AN22X2

MACRO AN22X1
    CLASS CORE ;
    FOREIGN AN22X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.959  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.055 2.895 3.030 3.235 ;
        RECT  2.800 1.010 3.030 3.235 ;
        RECT  2.625 1.010 3.030 1.410 ;
        RECT  1.370 1.010 3.030 1.350 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.580 1.500 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.090 2.250 1.920 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.945 1.640 2.570 2.020 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.424  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.190 0.600 2.630 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.760 3.540 1.100 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.565 -0.400 2.905 0.780 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.860 1.675 3.200 ;
        RECT  1.335 2.860 1.675 4.165 ;
        RECT  1.335 3.825 2.985 4.165 ;
    END
END AN22X1

MACRO AN22X0
    CLASS CORE ;
    FOREIGN AN22X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.849  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.310 2.310 2.650 3.660 ;
        RECT  2.170 1.010 2.400 2.540 ;
        RECT  1.995 1.010 2.400 1.410 ;
        RECT  1.370 1.010 2.400 1.350 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.153  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.560 1.270 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.153  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.220 1.940 2.630 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.153  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 1.530 3.035 2.080 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.153  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.195 0.600 2.775 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.740 3.930 1.080 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  2.630 -0.400 2.970 1.300 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 3.160 1.880 3.500 ;
        RECT  1.540 3.160 1.880 3.990 ;
    END
END AN22X0

MACRO AN222X4
    CLASS CORE ;
    FOREIGN AN222X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.895 2.195 4.475 2.635 ;
        RECT  3.995 2.120 4.475 2.635 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.295 1.610 3.825 1.950 ;
        RECT  3.295 1.610 3.665 2.635 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.375 2.230 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.605 1.915 2.220 2.255 ;
        RECT  1.605 1.030 1.870 2.255 ;
        RECT  1.385 1.030 1.870 1.410 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.490 2.120 3.065 2.635 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.961  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.510 2.920 8.010 3.260 ;
        RECT  6.400 1.360 8.010 1.700 ;
        RECT  7.055 1.360 7.435 3.260 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.020 0.515 1.590 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  7.090 3.560 7.430 5.280 ;
        RECT  5.855 3.555 6.195 5.280 ;
        RECT  1.620 3.840 1.960 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  7.035 -0.400 7.375 1.130 ;
        RECT  5.810 -0.400 6.150 1.090 ;
        RECT  3.330 -0.400 3.670 0.905 ;
        RECT  0.810 -0.400 1.150 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 3.325 2.700 3.555 ;
        RECT  0.900 3.325 1.240 4.180 ;
        RECT  2.360 3.325 2.700 4.180 ;
        RECT  0.180 2.865 3.420 3.095 ;
        RECT  3.080 2.865 3.420 4.160 ;
        RECT  0.180 2.865 0.520 4.160 ;
        RECT  4.520 3.345 4.860 4.160 ;
        RECT  3.080 3.840 4.860 4.160 ;
        RECT  4.520 1.025 4.935 1.365 ;
        RECT  2.100 1.135 4.935 1.365 ;
        RECT  2.100 0.880 2.440 1.685 ;
        RECT  4.705 2.120 5.115 2.460 ;
        RECT  4.705 1.025 4.935 3.095 ;
        RECT  3.800 2.865 4.935 3.095 ;
        RECT  3.800 2.865 4.140 3.450 ;
        RECT  5.220 1.360 5.575 1.700 ;
        RECT  5.345 1.945 6.500 2.285 ;
        RECT  5.345 1.360 5.575 3.260 ;
        RECT  5.220 2.915 5.575 3.260 ;
        RECT  0.180 2.865 2.30 3.095 ;
        RECT  2.100 1.135 3.40 1.365 ;
    END
END AN222X4

MACRO AN222X2
    CLASS CORE ;
    FOREIGN AN222X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.430 0.630 3.950 0.930 ;
        RECT  2.645 1.030 3.660 1.410 ;
        RECT  3.430 0.630 3.660 1.410 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.955 2.250 3.665 2.635 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.175 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.505 1.030 1.820 2.020 ;
        RECT  1.385 1.030 1.820 1.410 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.725 2.635 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.795 2.750 6.190 3.560 ;
        RECT  5.960 1.250 6.190 3.560 ;
        RECT  5.850 1.250 6.190 1.590 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.630 0.515 2.200 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  6.410 3.960 6.750 5.280 ;
        RECT  5.090 3.960 5.430 5.280 ;
        RECT  1.300 3.930 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  6.405 -0.400 6.750 0.720 ;
        RECT  5.285 -0.400 5.630 0.720 ;
        RECT  2.860 -0.400 3.200 0.710 ;
        RECT  0.555 -0.400 0.895 1.310 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 3.190 1.080 3.700 ;
        RECT  0.740 3.470 2.230 3.700 ;
        RECT  2.000 3.470 2.230 4.250 ;
        RECT  2.000 3.930 2.340 4.250 ;
        RECT  0.180 2.710 1.540 2.940 ;
        RECT  1.310 2.710 1.540 3.240 ;
        RECT  1.310 3.010 2.930 3.240 ;
        RECT  0.180 2.710 0.410 4.250 ;
        RECT  2.700 3.010 2.930 4.250 ;
        RECT  0.180 3.930 0.520 4.250 ;
        RECT  2.700 3.930 4.160 4.250 ;
        RECT  2.050 1.360 2.365 1.870 ;
        RECT  3.890 1.360 4.285 1.870 ;
        RECT  2.050 1.640 4.285 1.870 ;
        RECT  4.055 1.945 4.455 2.285 ;
        RECT  4.055 1.360 4.285 3.350 ;
        RECT  3.260 3.010 4.285 3.350 ;
        RECT  4.490 0.665 4.915 1.005 ;
        RECT  4.685 1.945 5.730 2.285 ;
        RECT  4.685 0.665 4.915 3.560 ;
        RECT  4.530 2.750 4.915 3.560 ;
        RECT  2.050 1.640 3.60 1.870 ;
    END
END AN222X2

MACRO AN222X1
    CLASS CORE ;
    FOREIGN AN222X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.525 1.480 4.915 2.170 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.295 2.120 3.825 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.375 2.230 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.430  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.605 1.915 2.220 2.255 ;
        RECT  1.605 1.030 1.870 2.255 ;
        RECT  1.385 1.030 1.870 1.410 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.490 2.120 3.065 2.635 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.903  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.055 0.910 4.860 1.250 ;
        RECT  3.800 2.860 4.285 3.450 ;
        RECT  4.055 0.910 4.285 3.450 ;
        RECT  2.100 1.455 4.285 1.685 ;
        RECT  2.100 0.880 2.440 1.685 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 0.980 0.515 1.590 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.040 5.280 ;
        RECT  1.620 3.840 1.960 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.040 0.400 ;
        RECT  3.330 -0.400 3.670 1.180 ;
        RECT  0.810 -0.400 1.150 1.410 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 3.325 2.700 3.555 ;
        RECT  0.900 3.325 1.240 4.180 ;
        RECT  2.360 3.325 2.700 4.180 ;
        RECT  0.180 2.865 3.420 3.095 ;
        RECT  3.080 2.865 3.420 4.160 ;
        RECT  0.180 2.865 0.520 4.160 ;
        RECT  4.520 2.865 4.860 4.160 ;
        RECT  3.080 3.840 4.860 4.160 ;
        RECT  0.180 2.865 2.50 3.095 ;
    END
END AN222X1

MACRO AN222X0
    CLASS CORE ;
    FOREIGN AN222X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN F
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.430 0.630 3.950 0.905 ;
        RECT  2.645 1.030 3.660 1.410 ;
        RECT  3.430 0.630 3.660 1.410 ;
        END
    END F
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.050 2.250 3.665 2.630 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.175 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.505 1.030 1.820 2.010 ;
        RECT  1.385 1.030 1.820 1.410 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 2.250 2.725 2.635 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.187  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.630 0.515 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.036  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.330 3.110 4.285 3.450 ;
        RECT  4.055 1.135 4.285 3.450 ;
        RECT  3.905 2.860 4.285 3.450 ;
        RECT  2.050 1.640 4.285 1.870 ;
        RECT  3.890 1.135 4.285 1.870 ;
        RECT  2.050 1.350 2.365 1.870 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.300 3.930 1.640 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  2.860 -0.400 3.200 0.710 ;
        RECT  0.555 -0.400 0.895 1.310 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.740 3.190 1.080 3.700 ;
        RECT  0.740 3.470 2.265 3.700 ;
        RECT  2.035 3.470 2.265 4.250 ;
        RECT  2.035 3.930 2.375 4.250 ;
        RECT  0.180 2.710 1.540 2.940 ;
        RECT  1.310 2.710 1.540 3.240 ;
        RECT  1.310 3.010 3.000 3.240 ;
        RECT  0.180 2.710 0.410 4.250 ;
        RECT  2.770 3.010 3.000 4.250 ;
        RECT  0.180 3.930 0.520 4.250 ;
        RECT  2.770 3.930 4.230 4.250 ;
    END
END AN222X0

MACRO AN221X4
    CLASS CORE ;
    FOREIGN AN221X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.190 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.840 2.170 4.235 2.630 ;
        RECT  3.615 2.170 4.235 2.460 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.640 1.525 2.220 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.955 3.385 2.295 ;
        RECT  2.625 1.640 3.045 2.295 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.905 1.640 2.395 2.220 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  7.670 0.890 8.010 3.560 ;
        RECT  6.230 2.250 8.010 2.630 ;
        RECT  6.230 0.890 6.570 3.560 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.010 0.510 1.640 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 8.190 5.280 ;
        RECT  6.950 2.860 7.290 5.280 ;
        RECT  5.510 2.750 5.850 5.280 ;
        RECT  1.675 3.610 2.015 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 8.190 0.400 ;
        RECT  6.950 -0.400 7.290 1.700 ;
        RECT  5.510 -0.400 5.850 1.700 ;
        RECT  3.325 -0.400 3.665 0.710 ;
        RECT  0.940 -0.400 1.280 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.905 3.150 2.775 3.380 ;
        RECT  0.905 3.150 1.245 4.065 ;
        RECT  2.435 3.150 2.775 4.065 ;
        RECT  0.180 2.690 3.610 2.920 ;
        RECT  0.180 2.690 0.520 4.180 ;
        RECT  3.270 2.690 3.610 4.180 ;
        RECT  2.135 0.975 4.425 1.340 ;
        RECT  4.195 0.975 4.425 1.940 ;
        RECT  4.195 1.710 4.630 1.940 ;
        RECT  4.465 1.945 4.750 2.285 ;
        RECT  4.465 1.775 4.695 3.090 ;
        RECT  4.050 2.860 4.695 3.090 ;
        RECT  4.050 2.860 4.415 4.205 ;
        RECT  4.790 0.780 5.210 1.540 ;
        RECT  4.980 1.945 6.000 2.285 ;
        RECT  4.980 0.780 5.210 4.180 ;
        RECT  4.785 3.370 5.210 4.180 ;
        RECT  0.180 2.690 2.20 2.920 ;
        RECT  2.135 0.975 3.60 1.340 ;
    END
END AN221X4

MACRO AN221X2
    CLASS CORE ;
    FOREIGN AN221X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.193  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.270 3.430 3.670 4.045 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.175 2.360 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.020 2.250 2.720 2.635 ;
        RECT  2.340 2.245 2.720 2.635 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.505 1.880 1.790 2.220 ;
        RECT  1.505 1.030 1.750 2.220 ;
        RECT  1.385 1.030 1.750 1.410 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.165 2.750 5.560 3.560 ;
        RECT  5.330 1.250 5.560 3.560 ;
        RECT  5.220 1.250 5.560 1.590 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.205  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 1.630 0.515 2.200 ;
        END
    END D
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.775 -0.400 6.120 0.720 ;
        RECT  4.655 -0.400 5.000 0.720 ;
        RECT  2.760 -0.400 3.100 0.960 ;
        RECT  0.500 -0.400 0.840 1.310 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 3.960 6.120 5.280 ;
        RECT  4.460 3.960 4.800 5.280 ;
        RECT  1.300 3.930 1.640 5.280 ;
        END
    END vdd!
    OBS
        LAYER MET1 ;
        RECT  0.740 3.190 1.080 3.700 ;
        RECT  0.740 3.470 2.230 3.700 ;
        RECT  2.000 3.470 2.230 4.250 ;
        RECT  2.000 3.930 2.340 4.250 ;
        RECT  0.180 2.730 1.540 2.960 ;
        RECT  1.310 2.730 1.540 3.240 ;
        RECT  1.310 3.010 2.930 3.240 ;
        RECT  0.180 2.730 0.410 4.250 ;
        RECT  2.700 3.010 2.930 4.250 ;
        RECT  0.180 3.930 0.520 4.250 ;
        RECT  2.700 3.930 3.040 4.250 ;
        RECT  1.980 1.360 3.700 1.700 ;
        RECT  3.425 1.360 3.700 2.285 ;
        RECT  3.425 1.945 3.850 2.285 ;
        RECT  3.425 1.360 3.655 2.980 ;
        RECT  3.300 2.640 3.655 2.980 ;
        RECT  3.860 0.665 4.310 1.005 ;
        RECT  4.080 1.945 5.100 2.285 ;
        RECT  4.080 0.665 4.310 3.560 ;
        RECT  3.900 3.220 4.310 3.560 ;
    END
END AN221X2

MACRO AN221X1
    CLASS CORE ;
    FOREIGN AN221X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.410 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.404  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.265 2.250 3.825 2.605 ;
        RECT  3.495 2.105 3.825 2.605 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.640 1.370 2.220 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.625 1.640 3.195 2.030 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.805 1.640 2.395 2.220 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.523  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.870 2.835 4.285 4.180 ;
        RECT  4.055 1.045 4.285 4.180 ;
        RECT  1.940 1.045 4.285 1.410 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.432  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 0.980 0.515 1.590 ;
        END
    END D
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 4.410 5.280 ;
        RECT  1.670 3.610 2.010 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 4.410 0.400 ;
        RECT  3.130 -0.400 3.470 0.815 ;
        RECT  0.790 -0.400 1.130 1.340 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.900 3.150 2.615 3.380 ;
        RECT  0.900 3.150 1.240 4.180 ;
        RECT  2.385 3.365 2.770 4.180 ;
        RECT  0.180 2.690 3.050 2.920 ;
        RECT  0.180 2.690 2.40 2.920 ;
        RECT  2.830 2.835 3.490 3.065 ;
        RECT  0.180 2.690 0.520 4.180 ;
        RECT  3.150 2.835 3.490 4.180 ;
    END
END AN221X1

MACRO AN221X0
    CLASS CORE ;
    FOREIGN AN221X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN E
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 2.300 3.205 2.760 ;
        END
    END E
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.740 1.640 1.155 2.455 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.015 1.640 2.765 2.070 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.690 2.300 2.030 2.585 ;
        RECT  1.385 2.030 1.785 2.580 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.182  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.030 0.505 2.085 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.195  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  3.260 3.470 3.665 4.250 ;
        RECT  3.435 0.630 3.665 4.250 ;
        RECT  1.475 1.180 3.665 1.410 ;
        RECT  3.260 0.630 3.665 1.410 ;
        RECT  1.475 0.630 1.815 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.340 3.930 1.680 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.505 -0.400 2.845 0.950 ;
        RECT  0.735 -0.400 1.075 0.970 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.760 3.270 1.100 3.680 ;
        RECT  0.760 3.450 2.380 3.680 ;
        RECT  2.040 3.450 2.380 4.250 ;
        RECT  0.290 2.810 1.560 3.040 ;
        RECT  1.330 2.990 3.030 3.220 ;
        RECT  2.700 2.990 3.030 3.440 ;
        RECT  0.290 2.810 0.520 4.250 ;
        RECT  0.180 3.930 0.520 4.250 ;
    END
END AN221X0

MACRO AN21X4
    CLASS CORE ;
    FOREIGN AN21X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.225 0.620 2.710 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.382  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.200 2.660 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.780 0.890 6.175 3.895 ;
        RECT  4.450 2.050 6.175 2.280 ;
        RECT  4.340 2.640 4.680 3.895 ;
        RECT  4.450 0.890 4.680 3.895 ;
        RECT  4.340 0.890 4.680 1.700 ;
        END
    END Q
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.400  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.510 2.020 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.060 2.640 5.400 5.280 ;
        RECT  3.620 2.640 3.960 5.280 ;
        RECT  0.900 3.400 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.060 -0.400 5.400 1.700 ;
        RECT  3.620 -0.400 3.960 1.700 ;
        RECT  2.200 -0.400 2.540 1.400 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.940 1.960 3.170 ;
        RECT  0.180 2.940 0.520 4.180 ;
        RECT  1.620 2.940 1.960 4.180 ;
        RECT  1.410 0.905 1.970 1.245 ;
        RECT  1.740 0.905 1.970 1.860 ;
        RECT  1.740 1.630 2.670 1.860 ;
        RECT  2.435 1.630 2.670 4.180 ;
        RECT  2.435 1.945 2.825 2.285 ;
        RECT  2.435 1.945 2.680 4.180 ;
        RECT  2.340 3.840 2.680 4.180 ;
        RECT  2.900 0.780 3.285 1.700 ;
        RECT  3.055 1.945 4.220 2.285 ;
        RECT  3.055 0.780 3.285 3.490 ;
        RECT  2.910 2.640 3.285 3.490 ;
    END
END AN21X4

MACRO AN21X2
    CLASS CORE ;
    FOREIGN AN21X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.825 2.250 2.420 2.660 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.525 2.020 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.200  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.220 0.640 2.660 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  4.430 2.880 4.915 3.690 ;
        RECT  4.535 0.950 4.915 3.690 ;
        RECT  4.430 0.950 4.915 1.290 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 5.670 5.280 ;
        RECT  5.150 2.815 5.490 5.280 ;
        RECT  3.670 4.090 4.010 5.280 ;
        RECT  0.900 3.350 1.240 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 5.670 0.400 ;
        RECT  5.150 -0.400 5.490 1.270 ;
        RECT  3.725 -0.400 4.050 1.270 ;
        RECT  2.215 -0.400 2.555 1.400 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.890 1.960 3.120 ;
        RECT  0.180 2.890 0.520 3.485 ;
        RECT  1.620 2.890 1.960 3.485 ;
        RECT  1.410 1.060 1.985 1.400 ;
        RECT  1.755 1.060 1.985 2.020 ;
        RECT  1.755 1.790 2.880 2.020 ;
        RECT  2.650 2.075 3.035 2.415 ;
        RECT  2.650 1.790 2.880 3.525 ;
        RECT  2.340 3.185 2.880 3.525 ;
        RECT  2.990 0.930 3.495 1.270 ;
        RECT  3.265 2.075 4.305 2.415 ;
        RECT  3.265 0.930 3.495 3.690 ;
        RECT  3.110 2.880 3.495 3.690 ;
    END
END AN21X2

MACRO AN21X1
    CLASS CORE ;
    FOREIGN AN21X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.026  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.935 2.450 2.275 4.105 ;
        RECT  1.605 2.450 2.275 2.680 ;
        RECT  1.605 1.030 1.835 2.680 ;
        RECT  1.330 1.030 1.835 1.420 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.120 1.635 0.525 2.395 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.413  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.065 1.505 2.405 2.220 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.434  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 2.240 1.375 2.635 ;
        END
    END A
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.755 3.790 1.095 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  2.000 -0.400 2.340 0.720 ;
        RECT  0.180 -0.400 0.520 1.400 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.985 1.670 3.325 ;
    END
END AN21X1

MACRO AN21X0
    CLASS CORE ;
    FOREIGN AN21X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.576  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.640 3.930 2.395 4.250 ;
        RECT  2.165 1.010 2.395 4.250 ;
        RECT  2.000 1.010 2.395 1.410 ;
        RECT  1.300 1.010 2.395 1.300 ;
        END
    END Q
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.158  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 1.030 0.525 1.990 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.158  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.530 1.355 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.151  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 1.935 2.630 ;
        RECT  1.650 1.735 1.935 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 2.520 5.280 ;
        RECT  0.880 3.650 1.220 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 2.520 0.400 ;
        RECT  2.000 -0.400 2.340 0.710 ;
        RECT  0.180 -0.400 0.520 0.710 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.955 1.935 3.295 ;
        RECT  0.180 2.955 0.520 3.990 ;
    END
END AN21X0

MACRO AN211X4
    CLASS CORE ;
    FOREIGN AN211X4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.417  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.420 2.175 2.975 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.080 0.525 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.470 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.269  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  6.410 0.890 6.750 3.560 ;
        RECT  4.970 2.250 6.750 2.630 ;
        RECT  4.970 0.890 5.310 3.560 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.417  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.190 2.630 ;
        RECT  1.850 2.175 2.190 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.930 5.280 ;
        RECT  5.690 2.860 6.030 5.280 ;
        RECT  4.250 2.750 4.590 5.280 ;
        RECT  0.940 3.370 1.280 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.930 0.400 ;
        RECT  5.690 -0.400 6.030 1.700 ;
        RECT  4.250 -0.400 4.590 1.700 ;
        RECT  2.160 -0.400 2.445 1.215 ;
        RECT  0.180 -0.400 0.520 1.490 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.860 2.000 3.140 ;
        RECT  0.180 2.860 0.520 4.140 ;
        RECT  1.660 2.860 2.000 4.170 ;
        RECT  1.370 0.885 1.930 1.225 ;
        RECT  1.700 0.885 1.930 1.945 ;
        RECT  2.810 0.885 3.165 1.945 ;
        RECT  1.700 1.715 3.385 1.945 ;
        RECT  3.205 1.765 3.525 2.285 ;
        RECT  3.205 1.765 3.445 3.090 ;
        RECT  2.810 2.860 3.445 3.090 ;
        RECT  2.810 2.860 3.150 4.170 ;
        RECT  3.530 0.780 3.985 1.535 ;
        RECT  3.755 1.945 4.740 2.285 ;
        RECT  3.755 0.780 3.985 4.180 ;
        RECT  3.530 3.320 3.985 4.180 ;
    END
END AN211X4

MACRO AN211X2
    CLASS CORE ;
    FOREIGN AN211X2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.206  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.460 2.120 2.985 2.630 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.222  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.120 0.545 2.630 ;
        RECT  0.115 1.915 0.525 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.222  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.470 2.020 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.896  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  5.060 2.860 5.545 3.560 ;
        RECT  5.060 1.250 5.400 3.560 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.206  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.230 2.630 ;
        RECT  1.850 2.010 2.230 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 6.300 5.280 ;
        RECT  5.780 2.750 6.120 5.280 ;
        RECT  4.340 2.750 4.680 5.280 ;
        RECT  0.980 3.430 1.320 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 6.300 0.400 ;
        RECT  5.780 -0.400 6.120 1.570 ;
        RECT  4.340 -0.400 4.680 1.570 ;
        RECT  2.170 -0.400 2.510 0.710 ;
        RECT  0.180 -0.400 0.520 1.310 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.180 2.860 2.080 3.200 ;
        RECT  1.370 1.070 3.230 1.410 ;
        RECT  3.000 1.070 3.230 1.890 ;
        RECT  3.215 1.945 3.605 2.285 ;
        RECT  3.215 1.660 3.445 3.230 ;
        RECT  2.890 2.890 3.445 3.230 ;
        RECT  3.580 1.120 4.065 1.460 ;
        RECT  3.835 1.945 4.830 2.285 ;
        RECT  3.835 1.120 4.065 3.560 ;
        RECT  3.675 2.750 4.065 3.560 ;
    END
END AN211X2

MACRO AN211X1
    CLASS CORE ;
    FOREIGN AN211X1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.417  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.645 1.640 3.175 2.160 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.125 2.120 0.625 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.448  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.170 1.640 1.715 2.035 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.542  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.890 2.640 3.655 3.260 ;
        RECT  3.405 1.070 3.655 3.260 ;
        RECT  1.450 1.070 3.655 1.410 ;
        RECT  2.890 2.640 3.230 4.170 ;
        END
    END Q
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.417  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.930 2.120 2.415 2.630 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.780 5.280 ;
        RECT  1.020 3.370 1.360 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.780 0.400 ;
        RECT  2.210 -0.400 2.550 0.840 ;
        RECT  0.260 -0.400 0.600 1.490 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.260 2.860 2.080 3.140 ;
        RECT  0.260 2.860 0.600 4.140 ;
        RECT  1.740 2.860 2.080 4.170 ;
    END
END AN211X1

MACRO AN211X0
    CLASS CORE ;
    FOREIGN AN211X0 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.150 BY 4.880 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.178  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.390 3.470 3.025 3.920 ;
        END
    END D
    PIN B
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.115 2.170 0.555 2.690 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.191  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  0.755 1.640 1.330 2.020 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAGATEAREA 0.178  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  1.385 2.250 2.060 2.630 ;
        RECT  1.720 2.025 2.060 2.630 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.842  LAYER MET1  ;
        PORT
        LAYER MET1 ;
        RECT  2.630 1.030 2.970 3.240 ;
        RECT  1.230 1.030 2.970 1.410 ;
        END
    END Q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 4.480 3.150 5.280 ;
        RECT  0.840 3.800 1.180 5.280 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER MET1 ;
        RECT  0.000 -0.400 3.150 0.400 ;
        RECT  1.930 -0.400 2.270 0.760 ;
        RECT  0.200 -0.400 0.540 0.760 ;
        END
    END gnd!
    OBS
        LAYER MET1 ;
        RECT  0.280 2.980 1.980 3.320 ;
        RECT  1.640 2.980 1.980 4.140 ;
    END
END AN211X0

END LIBRARY
