#************************************************************************/
# Copyright        : (c) All Rights Reserved
# Company          : X-FAB Semiconductor Foundries 
# Address          : Haarbergstr. 67,  D-99097 Erfurt, Germany
#
# File             : xc018_m6_FE.lef
# Description      : Layout Exchange Format
#                 
# Technology       : XC018M6
# Lib_version      : V 1.2.4
# Last Modified by : wad
# DATE             : Jul 11, 2007 
#
# Last Modified by : wad
# DATE             : Oct 19, 2007 
# descr            : new CAPACITANCE value
# DATE             : Jul  8, 2008
# desc             : add LOCKED layer
#
# DATE             : Sep  2, 2009
# desc             : add OVERLAP layer
#
# DATE             : Sep  28, 2009
# desc             : add INFLUENCE in wide metal rules
#
# DATE             : Sep 29, 2009 
# desc             : Modify VIARULE GENERATE
#************************************************************************/

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "<>" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID    0.005 ;
 
LAYER OVERLAP
   TYPE  OVERLAP ;
END OVERLAP

LAYER LOCKED
    TYPE MASTERSLICE ;
END LOCKED

LAYER LOCKED1
    TYPE MASTERSLICE ;
END LOCKED1

LAYER LOCKED2
    TYPE MASTERSLICE ;
END LOCKED2

LAYER MET1
    TYPE ROUTING ;
    WIDTH 0.230 ;
    SPACING 0.230 ;
    SPACING 0.600 RANGE 10.001 100 INFLUENCE 1.6 ;
    PITCH 0.610 ;
    OFFSET 0.000 ;
    AREA 0.202 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000076 ;
    EDGECAPACITANCE 0.000047 ;
    RESISTANCE RPERSQ 0.112 ;
    THICKNESS 0.62 ;
    ANTENNAAREARATIO 100 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFAREARATIO 9999999 ;
END MET1

LAYER VIA1
    TYPE CUT ;
END VIA1

LAYER MET2
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.600 RANGE 10.001 100 INFLUENCE 1.6 ;
    PITCH 0.630 ;
    OFFSET 0.315 ;
    AREA 0.202 ;
    WIREEXTENSION 0.19 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000081 ;
    EDGECAPACITANCE 0.000049 ;
    RESISTANCE RPERSQ 0.1 ;
    THICKNESS 0.62 ;
    ANTENNAAREARATIO 100 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFAREARATIO 9999999 ;
END MET2

LAYER VIA2
    TYPE CUT ;
END VIA2

LAYER MET3
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.600 RANGE 10.001 100 INFLUENCE 1.6 ;
    PITCH 0.610 ;
    OFFSET 0.000 ;
    AREA 0.202 ;
    WIREEXTENSION 0.19 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000081 ;
    EDGECAPACITANCE 0.000049 ;
    RESISTANCE RPERSQ 0.1 ;
    THICKNESS 0.62 ;
    ANTENNAAREARATIO 100 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFAREARATIO 9999999 ;
END MET3

LAYER VIA3
    TYPE CUT ;
END VIA3

LAYER MET4
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.600 RANGE 10.001 100 INFLUENCE 1.6 ;
    PITCH 0.630 ;
    OFFSET 0.315 ;
    AREA 0.202 ;
    WIREEXTENSION 0.19 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000081 ;
    EDGECAPACITANCE 0.000049 ;
    RESISTANCE RPERSQ 0.1 ;
    THICKNESS 0.62 ;
    ANTENNAAREARATIO 100 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFAREARATIO 9999999 ;
END MET4

LAYER VIA4
    TYPE CUT ;
END VIA4

LAYER MET5
    TYPE ROUTING ;
    WIDTH 0.280 ;
    SPACING 0.280 ;
    SPACING 0.600 RANGE 10.001 100 INFLUENCE 1.6 ;
    PITCH 0.610 ;
    OFFSET 0.000 ;
    AREA 0.202 ;
    WIREEXTENSION 0.19 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000075 ;
    EDGECAPACITANCE 0.000048 ;
    RESISTANCE RPERSQ 0.1 ;
    THICKNESS 0.62 ;
    ANTENNAAREARATIO 100 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFAREARATIO 9999999 ;
END MET5

LAYER VIATP
    TYPE CUT ;
END VIATP

LAYER METTP
    TYPE ROUTING ;
    WIDTH 0.440 ;
    SPACING 0.460 ;
    SPACING 0.600 RANGE 10.001 100 INFLUENCE 1.6 ;
    PITCH 1.260 ;
    OFFSET 0.315 ;
    AREA 0.562 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000034 ;
    EDGECAPACITANCE 0.000040 ;
    RESISTANCE RPERSQ 0.052 ;
    THICKNESS 1.09 ;
    ANTENNAAREARATIO 100 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFAREARATIO 9999999 ;
END METTP

VIA VIA1_X DEFAULT
    RESISTANCE 20.0 ;
    LAYER MET1 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA1 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET2 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA1_X

VIA VIA1_Y DEFAULT
    RESISTANCE 20.0 ;
    LAYER MET1 ;
        RECT -0.140 -0.190 0.140 0.190 ;
    LAYER VIA1 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET2 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA1_Y

VIA VIA2_small DEFAULT
    RESISTANCE 20.0 ;
    LAYER MET2 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA2_small

VIA VIA2_north DEFAULT TOPOFSTACKONLY
    RESISTANCE 20.0 ;
    LAYER MET2 ;
        RECT -0.140 -0.190 0.140 0.535 ;
    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA2_north

VIA VIA2_south DEFAULT TOPOFSTACKONLY
    RESISTANCE 20.0 ;
    LAYER MET2 ;
        RECT -0.140 -0.535 0.140 0.190 ;
    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA2_south

VIA VIA3_small DEFAULT
    RESISTANCE 20.0 ;
    LAYER MET3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA3_small

VIA VIA3_east DEFAULT TOPOFSTACKONLY
    RESISTANCE 20.0 ;
    LAYER MET3 ;
        RECT -0.190 -0.140 0.535 0.140 ;
    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA3_east

VIA VIA3_west DEFAULT TOPOFSTACKONLY
    RESISTANCE 20.0 ;
    LAYER MET3 ;
        RECT -0.535 -0.140 0.190 0.140 ;
    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA3_west

VIA VIA4_small DEFAULT
    RESISTANCE 20.0 ;
    LAYER MET4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET5 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA4_small

VIA VIA4_north DEFAULT TOPOFSTACKONLY
    RESISTANCE 20.0 ;
    LAYER MET4 ;
        RECT -0.140 -0.190 0.140 0.535 ;
    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET5 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA4_north

VIA VIA4_south DEFAULT TOPOFSTACKONLY
    RESISTANCE 20.0 ;
    LAYER MET4 ;
        RECT -0.140 -0.535 0.140 0.190 ;
    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER MET5 ;
        RECT -0.140 -0.140 0.140 0.140 ;
END VIA4_south

VIA VIATP_X DEFAULT
    RESISTANCE 13.0 ;
    LAYER MET5 ;
        RECT -0.270 -0.190 0.270 0.190 ;
    LAYER VIATP ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METTP ;
        RECT -0.270 -0.270 0.270 0.270 ;
END VIATP_X

VIA VIATP_Y DEFAULT
    RESISTANCE 13.0 ;
    LAYER MET5 ;
        RECT -0.190 -0.270 0.190 0.270 ;
    LAYER VIATP ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METTP ;
        RECT -0.270 -0.270 0.270 0.270 ;
END VIATP_Y

VIA VIA1_CH1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET1 ;
        RECT -0.190 -0.140 0.710 0.140 ;
    LAYER VIA1 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT  0.390 -0.130 0.650 0.130 ;
    LAYER MET2 ;
        RECT -0.140 -0.190 0.660 0.190 ;
END VIA1_CH1

VIA VIA1_CH2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET1 ;
        RECT -0.710 -0.140  0.190 0.140 ;
    LAYER VIA1 ;
        RECT -0.650 -0.130 -0.390 0.130 ;
        RECT -0.130 -0.130  0.130 0.130 ;
    LAYER MET2 ;
        RECT -0.660 -0.190  0.140 0.190 ;
END VIA1_CH2

VIA VIA1_CV1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET1 ;
        RECT -0.190 -0.660 0.190  0.140 ;
    LAYER VIA1 ;
        RECT -0.130 -0.130 0.130  0.130 ;
        RECT -0.130 -0.650 0.130 -0.390 ;
    LAYER MET2 ;
        RECT -0.140 -0.710 0.140  0.190 ;
END VIA1_CV1

VIA VIA1_CV2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET1 ;
        RECT -0.190 -0.140 0.190 0.660 ;
    LAYER VIA1 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT -0.130  0.390 0.130 0.650 ;
    LAYER MET2 ;
        RECT -0.140 -0.190 0.140 0.710 ;
END VIA1_CV2

VIA VIA2_CH1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET2 ;
        RECT -0.140 -0.190 0.660 0.190 ;
    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT  0.390 -0.130 0.650 0.130 ;
    LAYER MET3 ;
        RECT -0.190 -0.140 0.710 0.140 ;
END VIA2_CH1

VIA VIA2_CH2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET2 ;
        RECT -0.660 -0.190  0.140 0.190 ;
    LAYER VIA2 ;
        RECT -0.650 -0.130 -0.390 0.130 ;
        RECT -0.130 -0.130  0.130 0.130 ;
    LAYER MET3 ;
        RECT -0.710 -0.140  0.190 0.140 ;
END VIA2_CH2

VIA VIA2_CV1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET2 ;
        RECT -0.140 -0.710 0.140  0.190 ;
    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130  0.130 ;
        RECT -0.130 -0.650 0.130 -0.390 ;
    LAYER MET3 ;
        RECT -0.190 -0.660 0.190  0.140 ;
END VIA2_CV1

VIA VIA2_CV2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET2 ;
        RECT -0.140 -0.190 0.140 0.710 ;
    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT -0.130  0.390 0.130 0.650 ;
    LAYER MET3 ;
        RECT -0.190 -0.140 0.190 0.660 ;
END VIA2_CV2

VIA VIA3_CH1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET3 ;
        RECT -0.190 -0.140 0.710 0.140 ;
    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT  0.390 -0.130 0.650 0.130 ;
    LAYER MET4 ;
        RECT -0.140 -0.190 0.660 0.190 ;
END VIA3_CH1

VIA VIA3_CH2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET3 ;
        RECT -0.710 -0.140  0.190 0.140 ;
    LAYER VIA3 ;
        RECT -0.650 -0.130 -0.390 0.130 ;
        RECT -0.130 -0.130  0.130 0.130 ;
    LAYER MET4 ;
        RECT -0.660 -0.190  0.140 0.190 ;
END VIA3_CH2

VIA VIA3_CV1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET3 ;
        RECT -0.190 -0.660 0.190  0.140 ;
    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130  0.130 ;
        RECT -0.130 -0.650 0.130 -0.390 ;
    LAYER MET4 ;
        RECT -0.140 -0.710 0.140  0.190 ;
END VIA3_CV1

VIA VIA3_CV2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET3 ;
        RECT -0.190 -0.140 0.190 0.660 ;
    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT -0.130  0.390 0.130 0.650 ;
    LAYER MET4 ;
        RECT -0.140 -0.190 0.140 0.710 ;
END VIA3_CV2

VIA VIA4_CH1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET4 ;
        RECT -0.140 -0.190 0.660 0.190 ;
    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT  0.390 -0.130 0.650 0.130 ;
    LAYER MET5 ;
        RECT -0.190 -0.140 0.710 0.140 ;
END VIA4_CH1

VIA VIA4_CH2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET4 ;
        RECT -0.660 -0.190  0.140 0.190 ;
    LAYER VIA4 ;
        RECT -0.650 -0.130 -0.390 0.130 ;
        RECT -0.130 -0.130  0.130 0.130 ;
    LAYER MET5 ;
        RECT -0.710 -0.140  0.190 0.140 ;
END VIA4_CH2

VIA VIA4_CV1 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET4 ;
        RECT -0.140 -0.710 0.140  0.190 ;
    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130  0.130 ;
        RECT -0.130 -0.650 0.130 -0.390 ;
    LAYER MET5 ;
        RECT -0.190 -0.660 0.190  0.140 ;
END VIA4_CV1

VIA VIA4_CV2 DEFAULT
    RESISTANCE 10.0 ;
    LAYER MET4 ;
        RECT -0.140 -0.190 0.140 0.710 ;
    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        RECT -0.130  0.390 0.130 0.650 ;
    LAYER MET5 ;
        RECT -0.190 -0.140 0.190 0.660 ;
END VIA4_CV2

VIA VIATP_CH1 DEFAULT
    RESISTANCE 6.5 ;
    LAYER METTP ;
        RECT -0.270 -0.270 0.980 0.270 ;
    LAYER VIATP ;
        RECT -0.180 -0.180 0.180 0.180 ;
        RECT  0.530 -0.180 0.890 0.180 ;
    LAYER MET5 ;
        RECT -0.240 -0.190 0.950 0.190 ;
END VIATP_CH1

VIA VIATP_CH2 DEFAULT
    RESISTANCE 6.5 ;
    LAYER METTP ;
        RECT -0.980 -0.270  0.270 0.270 ;
    LAYER VIATP ;
        RECT -0.180 -0.180  0.180 0.180 ;
        RECT -0.890 -0.180 -0.530 0.180 ;
    LAYER MET5 ;
        RECT -0.950 -0.190  0.240 0.190 ;
END VIATP_CH2

VIA VIATP_CV1 DEFAULT
    RESISTANCE 6.5 ;
    LAYER METTP ;
        RECT -0.270 -0.980 0.270  0.270 ;
    LAYER VIATP ;
        RECT -0.180 -0.180 0.180  0.180 ;
        RECT -0.180 -0.890 0.180 -0.530 ;
    LAYER MET5 ;
        RECT -0.240 -0.900 0.240  0.190 ;
END VIATP_CV1

VIA VIATP_CV2 DEFAULT
    RESISTANCE 6.5 ;
    LAYER METTP ;
        RECT -0.270 -0.270 0.270 0.980 ;
    LAYER VIATP ;
        RECT -0.180 -0.180 0.180 0.180 ;
        RECT -0.180  0.530 0.180 0.890 ;
    LAYER MET5 ;
        RECT -0.240 -0.190 0.240 0.900 ;
END VIATP_CV2

VIARULE via1Array GENERATE
    LAYER MET1 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER MET2 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER VIA1 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
        RESISTANCE 20.0 ;
END via1Array

VIARULE via2Array GENERATE
    LAYER MET2 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER MET3 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER VIA2 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
        RESISTANCE 20.0 ;
END via2Array

VIARULE via3Array GENERATE
    LAYER MET3 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER MET4 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER VIA3 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
        RESISTANCE 20.0 ;
END via3Array

VIARULE via4Array GENERATE
    LAYER MET4 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER MET5 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER VIA4 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
        RESISTANCE 20.0 ;
END via4Array


VIARULE viaTPArray GENERATE
    LAYER MET5 ;
        ENCLOSURE 0.060 0.060 ;

    LAYER METTP ;
        ENCLOSURE 0.090 0.090 ;

    LAYER VIATP ;
        RECT -0.180 -0.180 0.180 0.180 ;
        SPACING 0.710 BY 0.710 ;
        RESISTANCE 13.0 ;
END viaTPArray

SPACING
    SAMENET MET1  MET1  0.230 STACK ;
    SAMENET MET2  MET2  0.280 STACK ;
    SAMENET MET3  MET3  0.280 STACK ;
    SAMENET MET4  MET4  0.280 STACK ;
    SAMENET MET5  MET5  0.280 STACK ;
    SAMENET METTP METTP 0.460 STACK ;
    SAMENET VIA1  VIA1  0.260 STACK ;
    SAMENET VIA2  VIA2  0.260 STACK ;
    SAMENET VIA3  VIA3  0.260 STACK ;
    SAMENET VIA4  VIA4  0.260 STACK ;
    SAMENET VIATP VIATP 0.350 STACK ;
    SAMENET VIA1  VIA2  0.0 STACK ;
    SAMENET VIA2  VIA3  0.0 STACK ;
    SAMENET VIA3  VIA4  0.0 STACK ;
    SAMENET VIA4  VIATP 0.0 STACK ;
END SPACING

END LIBRARY
